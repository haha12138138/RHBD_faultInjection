
module Custom_AES ( CLK, RSTn, EN, Kin, Din, KDrdy, Dout, Kvld, Dvld, BSY, 
        trigger );
  input [127:0] Kin;
  input [127:0] Din;
  output [127:0] Dout;
  input CLK, RSTn, EN, KDrdy;
  output Kvld, Dvld, BSY, trigger;
  wire [1:0] phase;
  wire   N0, KDrdy2, \U1/n1108 , \U1/n1107 , \U1/n1106 , \U1/n1105 ,
         \U1/n1104 , \U1/n1103 , \U1/n1102 , \U1/n1101 , \U1/n1100 ,
         \U1/n1099 , \U1/n1098 , \U1/n1097 , \U1/n1096 , \U1/n1095 , \U1/n670 ,
         \U1/n1 , \U1/n1094 , \U1/n1093 , \U1/n1092 , \U1/n1091 , \U1/n1090 ,
         \U1/n1089 , \U1/n1088 , \U1/n1087 , \U1/n1086 , \U1/n1085 ,
         \U1/n1084 , \U1/n1083 , \U1/n1082 , \U1/n1081 , \U1/n1080 ,
         \U1/n1079 , \U1/n1078 , \U1/n1077 , \U1/n1076 , \U1/n1075 ,
         \U1/n1074 , \U1/n1073 , \U1/n1072 , \U1/n1071 , \U1/n1070 ,
         \U1/n1069 , \U1/n1068 , \U1/n1067 , \U1/n1066 , \U1/n1065 ,
         \U1/n1064 , \U1/n1063 , \U1/n1062 , \U1/n1061 , \U1/n1060 ,
         \U1/n1059 , \U1/n1058 , \U1/n1057 , \U1/n1056 , \U1/n1055 ,
         \U1/n1054 , \U1/n1053 , \U1/n1052 , \U1/n1051 , \U1/n1050 ,
         \U1/n1049 , \U1/n1048 , \U1/n1047 , \U1/n1046 , \U1/n1045 ,
         \U1/n1044 , \U1/n1043 , \U1/n1042 , \U1/n1041 , \U1/n1040 ,
         \U1/n1039 , \U1/n1038 , \U1/n1037 , \U1/n1036 , \U1/n1035 ,
         \U1/n1034 , \U1/n1033 , \U1/n1032 , \U1/n1031 , \U1/n1030 ,
         \U1/n1029 , \U1/n1028 , \U1/n1027 , \U1/n1026 , \U1/n1025 ,
         \U1/n1024 , \U1/n1023 , \U1/n1022 , \U1/n1021 , \U1/n1020 ,
         \U1/n1019 , \U1/n1018 , \U1/n1017 , \U1/n1016 , \U1/n1015 ,
         \U1/n1014 , \U1/n1013 , \U1/n1012 , \U1/n1011 , \U1/n1010 ,
         \U1/n1009 , \U1/n1008 , \U1/n1007 , \U1/n1006 , \U1/n1005 ,
         \U1/n1004 , \U1/n1003 , \U1/n1002 , \U1/n1001 , \U1/n1000 , \U1/n999 ,
         \U1/n998 , \U1/n997 , \U1/n996 , \U1/n995 , \U1/n994 , \U1/n993 ,
         \U1/n992 , \U1/n991 , \U1/n990 , \U1/n989 , \U1/n988 , \U1/n987 ,
         \U1/n986 , \U1/n985 , \U1/n984 , \U1/n983 , \U1/n982 , \U1/n981 ,
         \U1/n980 , \U1/n979 , \U1/n978 , \U1/n977 , \U1/n976 , \U1/n975 ,
         \U1/n974 , \U1/n973 , \U1/n972 , \U1/n971 , \U1/n970 , \U1/n969 ,
         \U1/n968 , \U1/n967 , \U1/n966 , \U1/n965 , \U1/n964 , \U1/n963 ,
         \U1/n962 , \U1/n961 , \U1/n960 , \U1/n959 , \U1/n958 , \U1/n957 ,
         \U1/n956 , \U1/n955 , \U1/n954 , \U1/n953 , \U1/n952 , \U1/n951 ,
         \U1/n950 , \U1/n949 , \U1/n948 , \U1/n947 , \U1/n946 , \U1/n945 ,
         \U1/n944 , \U1/n943 , \U1/n942 , \U1/n941 , \U1/n940 , \U1/n939 ,
         \U1/n938 , \U1/n937 , \U1/n936 , \U1/n935 , \U1/n934 , \U1/n933 ,
         \U1/n932 , \U1/n931 , \U1/n930 , \U1/n929 , \U1/n928 , \U1/n927 ,
         \U1/n926 , \U1/n925 , \U1/n924 , \U1/n923 , \U1/n922 , \U1/n921 ,
         \U1/n920 , \U1/n919 , \U1/n918 , \U1/n917 , \U1/n916 , \U1/n915 ,
         \U1/n914 , \U1/n913 , \U1/n912 , \U1/n911 , \U1/n910 , \U1/n909 ,
         \U1/n908 , \U1/n907 , \U1/n906 , \U1/n905 , \U1/n904 , \U1/n903 ,
         \U1/n902 , \U1/n901 , \U1/n900 , \U1/n899 , \U1/n898 , \U1/n897 ,
         \U1/n896 , \U1/n895 , \U1/n894 , \U1/n893 , \U1/n892 , \U1/n891 ,
         \U1/n890 , \U1/n889 , \U1/n888 , \U1/n887 , \U1/n886 , \U1/n885 ,
         \U1/n884 , \U1/n883 , \U1/n882 , \U1/n881 , \U1/n880 , \U1/n879 ,
         \U1/n878 , \U1/n877 , \U1/n876 , \U1/n875 , \U1/n874 , \U1/n873 ,
         \U1/n872 , \U1/n871 , \U1/n870 , \U1/n869 , \U1/n868 , \U1/n867 ,
         \U1/n866 , \U1/n865 , \U1/n864 , \U1/n863 , \U1/n862 , \U1/n861 ,
         \U1/n860 , \U1/n859 , \U1/n858 , \U1/n857 , \U1/n856 , \U1/n855 ,
         \U1/n854 , \U1/n853 , \U1/n852 , \U1/n851 , \U1/n850 , \U1/n849 ,
         \U1/n848 , \U1/n847 , \U1/n846 , \U1/n845 , \U1/n844 , \U1/n843 ,
         \U1/n842 , \U1/n841 , \U1/n840 , \U1/n839 , \U1/n838 , \U1/n837 ,
         \U1/n836 , \U1/n835 , \U1/n834 , \U1/n833 , \U1/n832 , \U1/n831 ,
         \U1/n830 , \U1/n829 , \U1/n828 , \U1/n827 , \U1/n826 , \U1/n825 ,
         \U1/n824 , \U1/n823 , \U1/n822 , \U1/n821 , \U1/n820 , \U1/n819 ,
         \U1/n818 , \U1/n817 , \U1/n816 , \U1/n815 , \U1/n814 , \U1/n813 ,
         \U1/n812 , \U1/n811 , \U1/n810 , \U1/n809 , \U1/n808 , \U1/n807 ,
         \U1/n806 , \U1/n805 , \U1/n804 , \U1/n803 , \U1/n802 , \U1/n801 ,
         \U1/n800 , \U1/n799 , \U1/n798 , \U1/n797 , \U1/n796 , \U1/n795 ,
         \U1/n794 , \U1/n793 , \U1/n792 , \U1/n791 , \U1/n790 , \U1/n789 ,
         \U1/n788 , \U1/n787 , \U1/n786 , \U1/n785 , \U1/n784 , \U1/n783 ,
         \U1/n782 , \U1/n781 , \U1/n780 , \U1/n779 , \U1/n778 , \U1/n777 ,
         \U1/n776 , \U1/n775 , \U1/n774 , \U1/n773 , \U1/n772 , \U1/n771 ,
         \U1/n770 , \U1/n769 , \U1/n768 , \U1/n767 , \U1/n766 , \U1/n765 ,
         \U1/n764 , \U1/n763 , \U1/n762 , \U1/n761 , \U1/n760 , \U1/n759 ,
         \U1/n758 , \U1/n757 , \U1/n756 , \U1/n755 , \U1/n754 , \U1/n753 ,
         \U1/n752 , \U1/n751 , \U1/n750 , \U1/n749 , \U1/n748 , \U1/n747 ,
         \U1/n746 , \U1/n745 , \U1/n744 , \U1/n743 , \U1/n742 , \U1/n741 ,
         \U1/n740 , \U1/n739 , \U1/n738 , \U1/n737 , \U1/n736 , \U1/n735 ,
         \U1/n734 , \U1/n733 , \U1/n732 , \U1/n731 , \U1/n730 , \U1/n729 ,
         \U1/n728 , \U1/n727 , \U1/n726 , \U1/n725 , \U1/n724 , \U1/n723 ,
         \U1/n722 , \U1/n721 , \U1/n720 , \U1/n719 , \U1/n718 , \U1/n717 ,
         \U1/n716 , \U1/n715 , \U1/n714 , \U1/n713 , \U1/n712 , \U1/n711 ,
         \U1/n710 , \U1/n709 , \U1/n708 , \U1/n707 , \U1/n706 , \U1/n705 ,
         \U1/n704 , \U1/n703 , \U1/n702 , \U1/n701 , \U1/n700 , \U1/n699 ,
         \U1/n698 , \U1/n697 , \U1/n696 , \U1/n695 , \U1/n694 , \U1/n693 ,
         \U1/n692 , \U1/n691 , \U1/n690 , \U1/n689 , \U1/n688 , \U1/n687 ,
         \U1/n686 , \U1/n685 , \U1/n684 , \U1/n683 , \U1/n682 , \U1/n681 ,
         \U1/n680 , \U1/n679 , \U1/n678 , \U1/n677 , \U1/n676 , \U1/n675 ,
         \U1/n674 , \U1/n673 , \U1/n672 , \U1/n671 , \U1/n669 , \U1/n668 ,
         \U1/n667 , \U1/n666 , \U1/n665 , \U1/n664 , \U1/n663 , \U1/n662 ,
         \U1/n661 , \U1/n660 , \U1/n659 , \U1/n658 , \U1/n657 , \U1/n656 ,
         \U1/n655 , \U1/n654 , \U1/n653 , \U1/n652 , \U1/n651 , \U1/n650 ,
         \U1/n649 , \U1/n648 , \U1/n647 , \U1/n646 , \U1/n645 , \U1/n644 ,
         \U1/n643 , \U1/n642 , \U1/n641 , \U1/n640 , \U1/n639 , \U1/n638 ,
         \U1/n637 , \U1/n636 , \U1/n635 , \U1/n634 , \U1/n633 , \U1/n632 ,
         \U1/n631 , \U1/n630 , \U1/n629 , \U1/n628 , \U1/n627 , \U1/n626 ,
         \U1/n625 , \U1/n624 , \U1/n623 , \U1/n622 , \U1/n621 , \U1/n620 ,
         \U1/n619 , \U1/n618 , \U1/n617 , \U1/n616 , \U1/n615 , \U1/n614 ,
         \U1/n613 , \U1/n612 , \U1/n611 , \U1/n610 , \U1/n609 , \U1/n608 ,
         \U1/n607 , \U1/n606 , \U1/n605 , \U1/n604 , \U1/n603 , \U1/n602 ,
         \U1/n601 , \U1/n600 , \U1/n599 , \U1/n598 , \U1/n597 , \U1/n596 ,
         \U1/n595 , \U1/n594 , \U1/n593 , \U1/n592 , \U1/n591 , \U1/n590 ,
         \U1/n589 , \U1/n588 , \U1/n587 , \U1/n586 , \U1/n585 , \U1/n584 ,
         \U1/n583 , \U1/n582 , \U1/n581 , \U1/n580 , \U1/n579 , \U1/n578 ,
         \U1/n577 , \U1/n576 , \U1/n575 , \U1/n574 , \U1/n573 , \U1/n572 ,
         \U1/n571 , \U1/n570 , \U1/n569 , \U1/n568 , \U1/n567 , \U1/n566 ,
         \U1/n565 , \U1/n564 , \U1/n563 , \U1/n562 , \U1/n561 , \U1/n560 ,
         \U1/n559 , \U1/n558 , \U1/n557 , \U1/n556 , \U1/n555 , \U1/n554 ,
         \U1/n553 , \U1/n552 , \U1/n551 , \U1/n550 , \U1/n549 , \U1/n548 ,
         \U1/n547 , \U1/n546 , \U1/n545 , \U1/n544 , \U1/n543 , \U1/n542 ,
         \U1/n541 , \U1/n540 , \U1/n539 , \U1/n538 , \U1/n537 , \U1/n536 ,
         \U1/n535 , \U1/n534 , \U1/n533 , \U1/n532 , \U1/n531 , \U1/n530 ,
         \U1/n529 , \U1/n528 , \U1/n527 , \U1/n526 , \U1/n525 , \U1/n524 ,
         \U1/n523 , \U1/n522 , \U1/n521 , \U1/n520 , \U1/n519 , \U1/n518 ,
         \U1/n517 , \U1/n516 , \U1/n515 , \U1/n514 , \U1/n513 , \U1/n512 ,
         \U1/n511 , \U1/n510 , \U1/n509 , \U1/n508 , \U1/n507 , \U1/n506 ,
         \U1/n505 , \U1/n504 , \U1/n503 , \U1/n502 , \U1/n501 , \U1/n500 ,
         \U1/n499 , \U1/n498 , \U1/n497 , \U1/n496 , \U1/n495 , \U1/n494 ,
         \U1/n493 , \U1/n492 , \U1/n491 , \U1/n490 , \U1/n489 , \U1/n488 ,
         \U1/n487 , \U1/n486 , \U1/n485 , \U1/n484 , \U1/n483 , \U1/n482 ,
         \U1/n481 , \U1/n480 , \U1/n479 , \U1/n478 , \U1/n477 , \U1/n476 ,
         \U1/n475 , \U1/n474 , \U1/n473 , \U1/n472 , \U1/n471 , \U1/n470 ,
         \U1/n469 , \U1/n468 , \U1/n467 , \U1/n466 , \U1/n465 , \U1/n464 ,
         \U1/n463 , \U1/n462 , \U1/n461 , \U1/n460 , \U1/n459 , \U1/n458 ,
         \U1/n457 , \U1/n456 , \U1/n455 , \U1/n454 , \U1/n453 , \U1/n452 ,
         \U1/n451 , \U1/n450 , \U1/n449 , \U1/n448 , \U1/n447 , \U1/n446 ,
         \U1/n445 , \U1/n444 , \U1/n443 , \U1/n442 , \U1/n441 , \U1/n440 ,
         \U1/n439 , \U1/n438 , \U1/n437 , \U1/n436 , \U1/n435 , \U1/n434 ,
         \U1/n433 , \U1/n432 , \U1/n431 , \U1/n430 , \U1/n429 , \U1/n428 ,
         \U1/n427 , \U1/n426 , \U1/n425 , \U1/n424 , \U1/n423 , \U1/n422 ,
         \U1/n421 , \U1/n420 , \U1/n419 , \U1/n418 , \U1/n417 , \U1/n416 ,
         \U1/n415 , \U1/n414 , \U1/n413 , \U1/n412 , \U1/n411 , \U1/n410 ,
         \U1/n409 , \U1/n408 , \U1/n407 , \U1/n406 , \U1/n405 , \U1/n404 ,
         \U1/n403 , \U1/n402 , \U1/n401 , \U1/n400 , \U1/n399 , \U1/n398 ,
         \U1/n397 , \U1/n396 , \U1/n395 , \U1/n394 , \U1/n393 , \U1/n392 ,
         \U1/n391 , \U1/n390 , \U1/n389 , \U1/n388 , \U1/n387 , \U1/n386 ,
         \U1/n385 , \U1/n384 , \U1/n383 , \U1/n382 , \U1/n381 , \U1/n380 ,
         \U1/n379 , \U1/n378 , \U1/n377 , \U1/n376 , \U1/n375 , \U1/n374 ,
         \U1/n373 , \U1/n372 , \U1/n371 , \U1/n370 , \U1/n369 , \U1/n368 ,
         \U1/n367 , \U1/n366 , \U1/n365 , \U1/n364 , \U1/n363 , \U1/n362 ,
         \U1/n361 , \U1/n360 , \U1/n359 , \U1/n358 , \U1/n357 , \U1/n356 ,
         \U1/n355 , \U1/n354 , \U1/n353 , \U1/n352 , \U1/n351 , \U1/n350 ,
         \U1/n349 , \U1/n348 , \U1/n347 , \U1/n346 , \U1/n345 , \U1/n344 ,
         \U1/n343 , \U1/n342 , \U1/n341 , \U1/n340 , \U1/n339 , \U1/n338 ,
         \U1/n337 , \U1/n336 , \U1/n335 , \U1/n334 , \U1/n333 , \U1/n332 ,
         \U1/n331 , \U1/n330 , \U1/n329 , \U1/n328 , \U1/n327 , \U1/n326 ,
         \U1/n325 , \U1/n324 , \U1/n323 , \U1/n322 , \U1/n321 , \U1/n320 ,
         \U1/n319 , \U1/n318 , \U1/n317 , \U1/n316 , \U1/n315 , \U1/n314 ,
         \U1/n313 , \U1/n312 , \U1/n311 , \U1/n310 , \U1/n309 , \U1/n308 ,
         \U1/n307 , \U1/n306 , \U1/n305 , \U1/n304 , \U1/n303 , \U1/n302 ,
         \U1/n301 , \U1/n300 , \U1/n299 , \U1/n298 , \U1/n297 , \U1/n296 ,
         \U1/n295 , \U1/n294 , \U1/n293 , \U1/n292 , \U1/n291 , \U1/n290 ,
         \U1/n289 , \U1/n288 , \U1/n287 , \U1/n286 , \U1/n285 , \U1/n284 ,
         \U1/n283 , \U1/n282 , \U1/n281 , \U1/n280 , \U1/n279 , \U1/n278 ,
         \U1/n277 , \U1/n276 , \U1/n275 , \U1/n274 , \U1/n273 , \U1/n272 ,
         \U1/n271 , \U1/n270 , \U1/n269 , \U1/n268 , \U1/n267 , \U1/n266 ,
         \U1/n265 , \U1/n264 , \U1/n263 , \U1/n262 , \U1/n261 , \U1/n260 ,
         \U1/n259 , \U1/n258 , \U1/n257 , \U1/n256 , \U1/n255 , \U1/n254 ,
         \U1/n253 , \U1/n252 , \U1/n251 , \U1/n250 , \U1/n249 , \U1/n248 ,
         \U1/n247 , \U1/n246 , \U1/n245 , \U1/n244 , \U1/n243 , \U1/n242 ,
         \U1/n241 , \U1/n240 , \U1/n239 , \U1/n238 , \U1/n237 , \U1/n236 ,
         \U1/n235 , \U1/n234 , \U1/n233 , \U1/n232 , \U1/n231 , \U1/n230 ,
         \U1/n229 , \U1/n228 , \U1/n227 , \U1/n226 , \U1/n225 , \U1/n224 ,
         \U1/n223 , \U1/n222 , \U1/n221 , \U1/n220 , \U1/n219 , \U1/n218 ,
         \U1/n217 , \U1/n216 , \U1/n215 , \U1/n214 , \U1/n213 , \U1/n212 ,
         \U1/n211 , \U1/n210 , \U1/n209 , \U1/n208 , \U1/n207 , \U1/n206 ,
         \U1/n205 , \U1/n204 , \U1/n203 , \U1/n202 , \U1/n201 , \U1/n200 ,
         \U1/n199 , \U1/n198 , \U1/n197 , \U1/n196 , \U1/n195 , \U1/n194 ,
         \U1/n193 , \U1/n192 , \U1/n191 , \U1/n190 , \U1/n189 , \U1/n188 ,
         \U1/n187 , \U1/n186 , \U1/n185 , \U1/n184 , \U1/n183 , \U1/n182 ,
         \U1/n181 , \U1/n180 , \U1/n179 , \U1/n178 , \U1/n177 , \U1/n176 ,
         \U1/n175 , \U1/n174 , \U1/n173 , \U1/n172 , \U1/n171 , \U1/n170 ,
         \U1/n169 , \U1/n168 , \U1/n167 , \U1/n166 , \U1/n165 , \U1/n164 ,
         \U1/n163 , \U1/n162 , \U1/n161 , \U1/n160 , \U1/n159 , \U1/n158 ,
         \U1/n157 , \U1/n156 , \U1/n155 , \U1/n154 , \U1/n153 , \U1/n152 ,
         \U1/n151 , \U1/n150 , \U1/n149 , \U1/n148 , \U1/n147 , \U1/n146 ,
         \U1/n145 , \U1/n144 , \U1/n143 , \U1/n142 , \U1/n141 , \U1/n140 ,
         \U1/n139 , \U1/n138 , \U1/n137 , \U1/n136 , \U1/n135 , \U1/n134 ,
         \U1/n133 , \U1/n132 , \U1/n131 , \U1/n130 , \U1/n129 , \U1/n128 ,
         \U1/n127 , \U1/n126 , \U1/n125 , \U1/n124 , \U1/n123 , \U1/n122 ,
         \U1/n121 , \U1/n120 , \U1/n119 , \U1/n118 , \U1/n117 , \U1/n116 ,
         \U1/n115 , \U1/n114 , \U1/n113 , \U1/n112 , \U1/n111 , \U1/n110 ,
         \U1/n109 , \U1/n108 , \U1/n107 , \U1/n106 , \U1/n105 , \U1/n104 ,
         \U1/n103 , \U1/n102 , \U1/n101 , \U1/n100 , \U1/n99 , \U1/n98 ,
         \U1/n97 , \U1/n96 , \U1/n95 , \U1/n94 , \U1/n93 , \U1/n92 , \U1/n91 ,
         \U1/n90 , \U1/n89 , \U1/n88 , \U1/n87 , \U1/n86 , \U1/n85 , \U1/n84 ,
         \U1/n83 , \U1/n82 , \U1/n81 , \U1/n80 , \U1/n79 , \U1/n78 , \U1/n77 ,
         \U1/n76 , \U1/n75 , \U1/n74 , \U1/n73 , \U1/n72 , \U1/n71 , \U1/n70 ,
         \U1/n69 , \U1/n68 , \U1/n67 , \U1/n66 , \U1/n65 , \U1/n64 , \U1/n63 ,
         \U1/n62 , \U1/n61 , \U1/n60 , \U1/n59 , \U1/n58 , \U1/n57 , \U1/n56 ,
         \U1/n55 , \U1/n54 , \U1/n53 , \U1/n52 , \U1/n51 , \U1/n50 , \U1/n49 ,
         \U1/n48 , \U1/n47 , \U1/n46 , \U1/n45 , \U1/n44 , \U1/n43 , \U1/n42 ,
         \U1/n41 , \U1/n40 , \U1/n39 , \U1/n38 , \U1/n37 , \U1/n36 , \U1/n35 ,
         \U1/n34 , \U1/n33 , \U1/n32 , \U1/n31 , \U1/n30 , \U1/n29 , \U1/n28 ,
         \U1/n27 , \U1/n26 , \U1/n25 , \U1/n24 , \U1/n23 , \U1/n22 , \U1/n21 ,
         \U1/n20 , \U1/n19 , \U1/n18 , \U1/n17 , \U1/n16 , \U1/n15 , \U1/n14 ,
         \U1/n13 , \U1/n12 , \U1/n11 , \U1/n10 , \U1/n9 , \U1/n8 , \U1/n7 ,
         \U1/n6 , \U1/n5 , \U1/n4 , \U1/n3 , \U1/n2 , \U1/sel , \U1/rst ,
         \U1/aes_core/n258 , \U1/aes_core/n257 , \U1/aes_core/n256 ,
         \U1/aes_core/n255 , \U1/aes_core/n254 , \U1/aes_core/n253 ,
         \U1/aes_core/n252 , \U1/aes_core/n251 , \U1/aes_core/n250 ,
         \U1/aes_core/n249 , \U1/aes_core/n248 , \U1/aes_core/n247 ,
         \U1/aes_core/n246 , \U1/aes_core/n245 , \U1/aes_core/n244 ,
         \U1/aes_core/n243 , \U1/aes_core/n242 , \U1/aes_core/n241 ,
         \U1/aes_core/n240 , \U1/aes_core/n239 , \U1/aes_core/n238 ,
         \U1/aes_core/n237 , \U1/aes_core/n236 , \U1/aes_core/n235 ,
         \U1/aes_core/n234 , \U1/aes_core/n233 , \U1/aes_core/n232 ,
         \U1/aes_core/n231 , \U1/aes_core/n230 , \U1/aes_core/n229 ,
         \U1/aes_core/n228 , \U1/aes_core/n227 , \U1/aes_core/n226 ,
         \U1/aes_core/n225 , \U1/aes_core/n224 , \U1/aes_core/n223 ,
         \U1/aes_core/n222 , \U1/aes_core/n221 , \U1/aes_core/n220 ,
         \U1/aes_core/n219 , \U1/aes_core/n218 , \U1/aes_core/n217 ,
         \U1/aes_core/n216 , \U1/aes_core/n215 , \U1/aes_core/n214 ,
         \U1/aes_core/n213 , \U1/aes_core/n212 , \U1/aes_core/n211 ,
         \U1/aes_core/n210 , \U1/aes_core/n209 , \U1/aes_core/n208 ,
         \U1/aes_core/n207 , \U1/aes_core/n206 , \U1/aes_core/n205 ,
         \U1/aes_core/n204 , \U1/aes_core/n203 , \U1/aes_core/n202 ,
         \U1/aes_core/n201 , \U1/aes_core/n200 , \U1/aes_core/n199 ,
         \U1/aes_core/n198 , \U1/aes_core/n197 , \U1/aes_core/n196 ,
         \U1/aes_core/n195 , \U1/aes_core/n194 , \U1/aes_core/n193 ,
         \U1/aes_core/n192 , \U1/aes_core/n191 , \U1/aes_core/n190 ,
         \U1/aes_core/n189 , \U1/aes_core/n188 , \U1/aes_core/n187 ,
         \U1/aes_core/n186 , \U1/aes_core/n185 , \U1/aes_core/n184 ,
         \U1/aes_core/n183 , \U1/aes_core/n182 , \U1/aes_core/n181 ,
         \U1/aes_core/n180 , \U1/aes_core/n179 , \U1/aes_core/n178 ,
         \U1/aes_core/n177 , \U1/aes_core/n176 , \U1/aes_core/n175 ,
         \U1/aes_core/n174 , \U1/aes_core/n173 , \U1/aes_core/n172 ,
         \U1/aes_core/n171 , \U1/aes_core/n170 , \U1/aes_core/n169 ,
         \U1/aes_core/n168 , \U1/aes_core/n167 , \U1/aes_core/n166 ,
         \U1/aes_core/n165 , \U1/aes_core/n164 , \U1/aes_core/n163 ,
         \U1/aes_core/n162 , \U1/aes_core/n161 , \U1/aes_core/n160 ,
         \U1/aes_core/n159 , \U1/aes_core/n158 , \U1/aes_core/n157 ,
         \U1/aes_core/n156 , \U1/aes_core/n155 , \U1/aes_core/n154 ,
         \U1/aes_core/n153 , \U1/aes_core/n152 , \U1/aes_core/n151 ,
         \U1/aes_core/n150 , \U1/aes_core/n149 , \U1/aes_core/n148 ,
         \U1/aes_core/n147 , \U1/aes_core/n146 , \U1/aes_core/n145 ,
         \U1/aes_core/n144 , \U1/aes_core/n143 , \U1/aes_core/n142 ,
         \U1/aes_core/n141 , \U1/aes_core/n140 , \U1/aes_core/n139 ,
         \U1/aes_core/n138 , \U1/aes_core/n137 , \U1/aes_core/n136 ,
         \U1/aes_core/n135 , \U1/aes_core/n134 , \U1/aes_core/n133 ,
         \U1/aes_core/n132 , \U1/aes_core/n131 , \U1/aes_core/n130 ,
         \U1/aes_core/n129 , \U1/aes_core/n128 , \U1/aes_core/n127 ,
         \U1/aes_core/n126 , \U1/aes_core/n125 , \U1/aes_core/n124 ,
         \U1/aes_core/n123 , \U1/aes_core/n122 , \U1/aes_core/n121 ,
         \U1/aes_core/n120 , \U1/aes_core/n119 , \U1/aes_core/n118 ,
         \U1/aes_core/n117 , \U1/aes_core/n116 , \U1/aes_core/n115 ,
         \U1/aes_core/n114 , \U1/aes_core/n113 , \U1/aes_core/n112 ,
         \U1/aes_core/n111 , \U1/aes_core/n110 , \U1/aes_core/n109 ,
         \U1/aes_core/n108 , \U1/aes_core/n107 , \U1/aes_core/n106 ,
         \U1/aes_core/n105 , \U1/aes_core/n104 , \U1/aes_core/n103 ,
         \U1/aes_core/n102 , \U1/aes_core/n101 , \U1/aes_core/n100 ,
         \U1/aes_core/n99 , \U1/aes_core/n98 , \U1/aes_core/n97 ,
         \U1/aes_core/n96 , \U1/aes_core/n95 , \U1/aes_core/n94 ,
         \U1/aes_core/n93 , \U1/aes_core/n92 , \U1/aes_core/n91 ,
         \U1/aes_core/n90 , \U1/aes_core/n89 , \U1/aes_core/n88 ,
         \U1/aes_core/n87 , \U1/aes_core/n86 , \U1/aes_core/n85 ,
         \U1/aes_core/n84 , \U1/aes_core/n83 , \U1/aes_core/n82 ,
         \U1/aes_core/n81 , \U1/aes_core/n80 , \U1/aes_core/n79 ,
         \U1/aes_core/n78 , \U1/aes_core/n77 , \U1/aes_core/n76 ,
         \U1/aes_core/n75 , \U1/aes_core/n74 , \U1/aes_core/n73 ,
         \U1/aes_core/n72 , \U1/aes_core/n71 , \U1/aes_core/n70 ,
         \U1/aes_core/n69 , \U1/aes_core/n68 , \U1/aes_core/n67 ,
         \U1/aes_core/n66 , \U1/aes_core/n65 , \U1/aes_core/n64 ,
         \U1/aes_core/n63 , \U1/aes_core/n62 , \U1/aes_core/n61 ,
         \U1/aes_core/n60 , \U1/aes_core/n59 , \U1/aes_core/n58 ,
         \U1/aes_core/n57 , \U1/aes_core/n56 , \U1/aes_core/n55 ,
         \U1/aes_core/n54 , \U1/aes_core/n53 , \U1/aes_core/n52 ,
         \U1/aes_core/n51 , \U1/aes_core/n50 , \U1/aes_core/n49 ,
         \U1/aes_core/n48 , \U1/aes_core/n47 , \U1/aes_core/n46 ,
         \U1/aes_core/n45 , \U1/aes_core/n44 , \U1/aes_core/n43 ,
         \U1/aes_core/n42 , \U1/aes_core/n41 , \U1/aes_core/n40 ,
         \U1/aes_core/n39 , \U1/aes_core/n38 , \U1/aes_core/n37 ,
         \U1/aes_core/n36 , \U1/aes_core/n35 , \U1/aes_core/n34 ,
         \U1/aes_core/n33 , \U1/aes_core/n32 , \U1/aes_core/n31 ,
         \U1/aes_core/n30 , \U1/aes_core/n29 , \U1/aes_core/n28 ,
         \U1/aes_core/n27 , \U1/aes_core/n26 , \U1/aes_core/n25 ,
         \U1/aes_core/n24 , \U1/aes_core/n23 , \U1/aes_core/n22 ,
         \U1/aes_core/n21 , \U1/aes_core/n20 , \U1/aes_core/n19 ,
         \U1/aes_core/n18 , \U1/aes_core/n17 , \U1/aes_core/n16 ,
         \U1/aes_core/n15 , \U1/aes_core/n14 , \U1/aes_core/n13 ,
         \U1/aes_core/n12 , \U1/aes_core/n11 , \U1/aes_core/n10 ,
         \U1/aes_core/n9 , \U1/aes_core/n8 , \U1/aes_core/n7 ,
         \U1/aes_core/n6 , \U1/aes_core/n5 , \U1/aes_core/n4 ,
         \U1/aes_core/n3 , \U1/aes_core/n2 , \U1/aes_core/n1 ,
         \U1/aes_core/SB0/n1690 , \U1/aes_core/SB0/n1689 ,
         \U1/aes_core/SB0/n1688 , \U1/aes_core/SB0/n1687 ,
         \U1/aes_core/SB0/n1686 , \U1/aes_core/SB0/n1685 ,
         \U1/aes_core/SB0/n1684 , \U1/aes_core/SB0/n1683 ,
         \U1/aes_core/SB0/n1682 , \U1/aes_core/SB0/n1681 ,
         \U1/aes_core/SB0/n1680 , \U1/aes_core/SB0/n1679 ,
         \U1/aes_core/SB0/n1678 , \U1/aes_core/SB0/n1677 ,
         \U1/aes_core/SB0/n1676 , \U1/aes_core/SB0/n1675 ,
         \U1/aes_core/SB0/n1674 , \U1/aes_core/SB0/n1673 ,
         \U1/aes_core/SB0/n1672 , \U1/aes_core/SB0/n1671 ,
         \U1/aes_core/SB0/n1670 , \U1/aes_core/SB0/n1669 ,
         \U1/aes_core/SB0/n1668 , \U1/aes_core/SB0/n1667 ,
         \U1/aes_core/SB0/n1666 , \U1/aes_core/SB0/n1665 ,
         \U1/aes_core/SB0/n1664 , \U1/aes_core/SB0/n1663 ,
         \U1/aes_core/SB0/n1662 , \U1/aes_core/SB0/n1661 ,
         \U1/aes_core/SB0/n1660 , \U1/aes_core/SB0/n1659 ,
         \U1/aes_core/SB0/n1658 , \U1/aes_core/SB0/n1657 ,
         \U1/aes_core/SB0/n1656 , \U1/aes_core/SB0/n1655 ,
         \U1/aes_core/SB0/n1654 , \U1/aes_core/SB0/n1653 ,
         \U1/aes_core/SB0/n1652 , \U1/aes_core/SB0/n1651 ,
         \U1/aes_core/SB0/n1650 , \U1/aes_core/SB0/n1649 ,
         \U1/aes_core/SB0/n1648 , \U1/aes_core/SB0/n1647 ,
         \U1/aes_core/SB0/n1646 , \U1/aes_core/SB0/n1645 ,
         \U1/aes_core/SB0/n1644 , \U1/aes_core/SB0/n1643 ,
         \U1/aes_core/SB0/n1642 , \U1/aes_core/SB0/n1641 ,
         \U1/aes_core/SB0/n1640 , \U1/aes_core/SB0/n1639 ,
         \U1/aes_core/SB0/n1638 , \U1/aes_core/SB0/n1637 ,
         \U1/aes_core/SB0/n1636 , \U1/aes_core/SB0/n1635 ,
         \U1/aes_core/SB0/n1634 , \U1/aes_core/SB0/n1633 ,
         \U1/aes_core/SB0/n1632 , \U1/aes_core/SB0/n1631 ,
         \U1/aes_core/SB0/n1630 , \U1/aes_core/SB0/n1629 ,
         \U1/aes_core/SB0/n1628 , \U1/aes_core/SB0/n1627 ,
         \U1/aes_core/SB0/n1626 , \U1/aes_core/SB0/n1625 ,
         \U1/aes_core/SB0/n1624 , \U1/aes_core/SB0/n1623 ,
         \U1/aes_core/SB0/n1622 , \U1/aes_core/SB0/n1620 ,
         \U1/aes_core/SB0/n1619 , \U1/aes_core/SB0/n1618 ,
         \U1/aes_core/SB0/n1617 , \U1/aes_core/SB0/n1616 ,
         \U1/aes_core/SB0/n1615 , \U1/aes_core/SB0/n1614 ,
         \U1/aes_core/SB0/n1613 , \U1/aes_core/SB0/n1612 ,
         \U1/aes_core/SB0/n1611 , \U1/aes_core/SB0/n1610 ,
         \U1/aes_core/SB0/n1609 , \U1/aes_core/SB0/n1608 ,
         \U1/aes_core/SB0/n1607 , \U1/aes_core/SB0/n1606 ,
         \U1/aes_core/SB0/n1605 , \U1/aes_core/SB0/n1604 ,
         \U1/aes_core/SB0/n1603 , \U1/aes_core/SB0/n1602 ,
         \U1/aes_core/SB0/n1601 , \U1/aes_core/SB0/n1600 ,
         \U1/aes_core/SB0/n1599 , \U1/aes_core/SB0/n1598 ,
         \U1/aes_core/SB0/n1597 , \U1/aes_core/SB0/n1596 ,
         \U1/aes_core/SB0/n1595 , \U1/aes_core/SB0/n1594 ,
         \U1/aes_core/SB0/n1593 , \U1/aes_core/SB0/n1592 ,
         \U1/aes_core/SB0/n1591 , \U1/aes_core/SB0/n1590 ,
         \U1/aes_core/SB0/n1589 , \U1/aes_core/SB0/n1588 ,
         \U1/aes_core/SB0/n1587 , \U1/aes_core/SB0/n1586 ,
         \U1/aes_core/SB0/n1585 , \U1/aes_core/SB0/n1584 ,
         \U1/aes_core/SB0/n1583 , \U1/aes_core/SB0/n1582 ,
         \U1/aes_core/SB0/n1581 , \U1/aes_core/SB0/n1580 ,
         \U1/aes_core/SB0/n1579 , \U1/aes_core/SB0/n1578 ,
         \U1/aes_core/SB0/n1577 , \U1/aes_core/SB0/n1576 ,
         \U1/aes_core/SB0/n1575 , \U1/aes_core/SB0/n1574 ,
         \U1/aes_core/SB0/n1573 , \U1/aes_core/SB0/n1572 ,
         \U1/aes_core/SB0/n1571 , \U1/aes_core/SB0/n1570 ,
         \U1/aes_core/SB0/n1569 , \U1/aes_core/SB0/n1568 ,
         \U1/aes_core/SB0/n1567 , \U1/aes_core/SB0/n1566 ,
         \U1/aes_core/SB0/n1565 , \U1/aes_core/SB0/n1564 ,
         \U1/aes_core/SB0/n1563 , \U1/aes_core/SB0/n1562 ,
         \U1/aes_core/SB0/n1561 , \U1/aes_core/SB0/n1560 ,
         \U1/aes_core/SB0/n1559 , \U1/aes_core/SB0/n1558 ,
         \U1/aes_core/SB0/n1557 , \U1/aes_core/SB0/n1556 ,
         \U1/aes_core/SB0/n1555 , \U1/aes_core/SB0/n1554 ,
         \U1/aes_core/SB0/n1553 , \U1/aes_core/SB0/n1552 ,
         \U1/aes_core/SB0/n1551 , \U1/aes_core/SB0/n1550 ,
         \U1/aes_core/SB0/n1549 , \U1/aes_core/SB0/n1548 ,
         \U1/aes_core/SB0/n1547 , \U1/aes_core/SB0/n1546 ,
         \U1/aes_core/SB0/n1545 , \U1/aes_core/SB0/n1544 ,
         \U1/aes_core/SB0/n1543 , \U1/aes_core/SB0/n1542 ,
         \U1/aes_core/SB0/n1541 , \U1/aes_core/SB0/n1540 ,
         \U1/aes_core/SB0/n1539 , \U1/aes_core/SB0/n1538 ,
         \U1/aes_core/SB0/n1537 , \U1/aes_core/SB0/n1536 ,
         \U1/aes_core/SB0/n1535 , \U1/aes_core/SB0/n1534 ,
         \U1/aes_core/SB0/n1533 , \U1/aes_core/SB0/n1532 ,
         \U1/aes_core/SB0/n1531 , \U1/aes_core/SB0/n1530 ,
         \U1/aes_core/SB0/n1529 , \U1/aes_core/SB0/n1528 ,
         \U1/aes_core/SB0/n1527 , \U1/aes_core/SB0/n1526 ,
         \U1/aes_core/SB0/n1525 , \U1/aes_core/SB0/n1524 ,
         \U1/aes_core/SB0/n1523 , \U1/aes_core/SB0/n1522 ,
         \U1/aes_core/SB0/n1521 , \U1/aes_core/SB0/n1520 ,
         \U1/aes_core/SB0/n1519 , \U1/aes_core/SB0/n1518 ,
         \U1/aes_core/SB0/n1517 , \U1/aes_core/SB0/n1516 ,
         \U1/aes_core/SB0/n1515 , \U1/aes_core/SB0/n1514 ,
         \U1/aes_core/SB0/n1513 , \U1/aes_core/SB0/n1512 ,
         \U1/aes_core/SB0/n1511 , \U1/aes_core/SB0/n1510 ,
         \U1/aes_core/SB0/n1509 , \U1/aes_core/SB0/n1508 ,
         \U1/aes_core/SB0/n1507 , \U1/aes_core/SB0/n1506 ,
         \U1/aes_core/SB0/n1505 , \U1/aes_core/SB0/n1504 ,
         \U1/aes_core/SB0/n1503 , \U1/aes_core/SB0/n1502 ,
         \U1/aes_core/SB0/n1501 , \U1/aes_core/SB0/n1500 ,
         \U1/aes_core/SB0/n1499 , \U1/aes_core/SB0/n1498 ,
         \U1/aes_core/SB0/n1497 , \U1/aes_core/SB0/n1496 ,
         \U1/aes_core/SB0/n1495 , \U1/aes_core/SB0/n1494 ,
         \U1/aes_core/SB0/n1493 , \U1/aes_core/SB0/n1492 ,
         \U1/aes_core/SB0/n1491 , \U1/aes_core/SB0/n1490 ,
         \U1/aes_core/SB0/n1489 , \U1/aes_core/SB0/n1488 ,
         \U1/aes_core/SB0/n1487 , \U1/aes_core/SB0/n1486 ,
         \U1/aes_core/SB0/n1485 , \U1/aes_core/SB0/n1484 ,
         \U1/aes_core/SB0/n1483 , \U1/aes_core/SB0/n1482 ,
         \U1/aes_core/SB0/n1481 , \U1/aes_core/SB0/n1480 ,
         \U1/aes_core/SB0/n1479 , \U1/aes_core/SB0/n1478 ,
         \U1/aes_core/SB0/n1477 , \U1/aes_core/SB0/n1476 ,
         \U1/aes_core/SB0/n1475 , \U1/aes_core/SB0/n1474 ,
         \U1/aes_core/SB0/n1473 , \U1/aes_core/SB0/n1472 ,
         \U1/aes_core/SB0/n1471 , \U1/aes_core/SB0/n1470 ,
         \U1/aes_core/SB0/n1469 , \U1/aes_core/SB0/n1468 ,
         \U1/aes_core/SB0/n1467 , \U1/aes_core/SB0/n1466 ,
         \U1/aes_core/SB0/n1465 , \U1/aes_core/SB0/n1464 ,
         \U1/aes_core/SB0/n1463 , \U1/aes_core/SB0/n1462 ,
         \U1/aes_core/SB0/n1461 , \U1/aes_core/SB0/n1460 ,
         \U1/aes_core/SB0/n1459 , \U1/aes_core/SB0/n1458 ,
         \U1/aes_core/SB0/n1457 , \U1/aes_core/SB0/n1456 ,
         \U1/aes_core/SB0/n1455 , \U1/aes_core/SB0/n1454 ,
         \U1/aes_core/SB0/n1453 , \U1/aes_core/SB0/n1452 ,
         \U1/aes_core/SB0/n1451 , \U1/aes_core/SB0/n1450 ,
         \U1/aes_core/SB0/n1449 , \U1/aes_core/SB0/n1448 ,
         \U1/aes_core/SB0/n1447 , \U1/aes_core/SB0/n1446 ,
         \U1/aes_core/SB0/n1445 , \U1/aes_core/SB0/n1444 ,
         \U1/aes_core/SB0/n1443 , \U1/aes_core/SB0/n1442 ,
         \U1/aes_core/SB0/n1441 , \U1/aes_core/SB0/n1440 ,
         \U1/aes_core/SB0/n1439 , \U1/aes_core/SB0/n1438 ,
         \U1/aes_core/SB0/n1437 , \U1/aes_core/SB0/n1436 ,
         \U1/aes_core/SB0/n1435 , \U1/aes_core/SB0/n1434 ,
         \U1/aes_core/SB0/n1433 , \U1/aes_core/SB0/n1432 ,
         \U1/aes_core/SB0/n1431 , \U1/aes_core/SB0/n1430 ,
         \U1/aes_core/SB0/n1429 , \U1/aes_core/SB0/n1428 ,
         \U1/aes_core/SB0/n1427 , \U1/aes_core/SB0/n1426 ,
         \U1/aes_core/SB0/n1425 , \U1/aes_core/SB0/n1424 ,
         \U1/aes_core/SB0/n1423 , \U1/aes_core/SB0/n1422 ,
         \U1/aes_core/SB0/n1421 , \U1/aes_core/SB0/n1420 ,
         \U1/aes_core/SB0/n1419 , \U1/aes_core/SB0/n1418 ,
         \U1/aes_core/SB0/n1417 , \U1/aes_core/SB0/n1416 ,
         \U1/aes_core/SB0/n1415 , \U1/aes_core/SB0/n1414 ,
         \U1/aes_core/SB0/n1413 , \U1/aes_core/SB0/n1412 ,
         \U1/aes_core/SB0/n1411 , \U1/aes_core/SB0/n1410 ,
         \U1/aes_core/SB0/n1409 , \U1/aes_core/SB0/n1408 ,
         \U1/aes_core/SB0/n1407 , \U1/aes_core/SB0/n1406 ,
         \U1/aes_core/SB0/n1405 , \U1/aes_core/SB0/n1404 ,
         \U1/aes_core/SB0/n1403 , \U1/aes_core/SB0/n1402 ,
         \U1/aes_core/SB0/n1401 , \U1/aes_core/SB0/n1400 ,
         \U1/aes_core/SB0/n1399 , \U1/aes_core/SB0/n1398 ,
         \U1/aes_core/SB0/n1397 , \U1/aes_core/SB0/n1396 ,
         \U1/aes_core/SB0/n1395 , \U1/aes_core/SB0/n1394 ,
         \U1/aes_core/SB0/n1393 , \U1/aes_core/SB0/n1392 ,
         \U1/aes_core/SB0/n1391 , \U1/aes_core/SB0/n1390 ,
         \U1/aes_core/SB0/n1389 , \U1/aes_core/SB0/n1388 ,
         \U1/aes_core/SB0/n1387 , \U1/aes_core/SB0/n1386 ,
         \U1/aes_core/SB0/n1385 , \U1/aes_core/SB0/n1384 ,
         \U1/aes_core/SB0/n1383 , \U1/aes_core/SB0/n1382 ,
         \U1/aes_core/SB0/n1381 , \U1/aes_core/SB0/n1380 ,
         \U1/aes_core/SB0/n1379 , \U1/aes_core/SB0/n1378 ,
         \U1/aes_core/SB0/n1377 , \U1/aes_core/SB0/n1376 ,
         \U1/aes_core/SB0/n1375 , \U1/aes_core/SB0/n1374 ,
         \U1/aes_core/SB0/n1373 , \U1/aes_core/SB0/n1372 ,
         \U1/aes_core/SB0/n1371 , \U1/aes_core/SB0/n1370 ,
         \U1/aes_core/SB0/n1369 , \U1/aes_core/SB0/n1368 ,
         \U1/aes_core/SB0/n1367 , \U1/aes_core/SB0/n1366 ,
         \U1/aes_core/SB0/n1365 , \U1/aes_core/SB0/n1364 ,
         \U1/aes_core/SB0/n1363 , \U1/aes_core/SB0/n1362 ,
         \U1/aes_core/SB0/n1361 , \U1/aes_core/SB0/n1360 ,
         \U1/aes_core/SB0/n1359 , \U1/aes_core/SB0/n1358 ,
         \U1/aes_core/SB0/n1357 , \U1/aes_core/SB0/n1356 ,
         \U1/aes_core/SB0/n1355 , \U1/aes_core/SB0/n1354 ,
         \U1/aes_core/SB0/n1353 , \U1/aes_core/SB0/n1352 ,
         \U1/aes_core/SB0/n1351 , \U1/aes_core/SB0/n1350 ,
         \U1/aes_core/SB0/n1349 , \U1/aes_core/SB0/n1348 ,
         \U1/aes_core/SB0/n1347 , \U1/aes_core/SB0/n1346 ,
         \U1/aes_core/SB0/n1345 , \U1/aes_core/SB0/n1344 ,
         \U1/aes_core/SB0/n1343 , \U1/aes_core/SB0/n1342 ,
         \U1/aes_core/SB0/n1341 , \U1/aes_core/SB0/n1340 ,
         \U1/aes_core/SB0/n1339 , \U1/aes_core/SB0/n1338 ,
         \U1/aes_core/SB0/n1337 , \U1/aes_core/SB0/n1336 ,
         \U1/aes_core/SB0/n1335 , \U1/aes_core/SB0/n1334 ,
         \U1/aes_core/SB0/n1333 , \U1/aes_core/SB0/n1332 ,
         \U1/aes_core/SB0/n1331 , \U1/aes_core/SB0/n1330 ,
         \U1/aes_core/SB0/n1329 , \U1/aes_core/SB0/n1328 ,
         \U1/aes_core/SB0/n1327 , \U1/aes_core/SB0/n1326 ,
         \U1/aes_core/SB0/n1325 , \U1/aes_core/SB0/n1324 ,
         \U1/aes_core/SB0/n1323 , \U1/aes_core/SB0/n1322 ,
         \U1/aes_core/SB0/n1321 , \U1/aes_core/SB0/n1320 ,
         \U1/aes_core/SB0/n1319 , \U1/aes_core/SB0/n1318 ,
         \U1/aes_core/SB0/n1317 , \U1/aes_core/SB0/n1316 ,
         \U1/aes_core/SB0/n1315 , \U1/aes_core/SB0/n1314 ,
         \U1/aes_core/SB0/n1313 , \U1/aes_core/SB0/n1312 ,
         \U1/aes_core/SB0/n1311 , \U1/aes_core/SB0/n1310 ,
         \U1/aes_core/SB0/n1309 , \U1/aes_core/SB0/n1308 ,
         \U1/aes_core/SB0/n1307 , \U1/aes_core/SB0/n1306 ,
         \U1/aes_core/SB0/n1305 , \U1/aes_core/SB0/n1304 ,
         \U1/aes_core/SB0/n1303 , \U1/aes_core/SB0/n1302 ,
         \U1/aes_core/SB0/n1301 , \U1/aes_core/SB0/n1300 ,
         \U1/aes_core/SB0/n1299 , \U1/aes_core/SB0/n1298 ,
         \U1/aes_core/SB0/n1297 , \U1/aes_core/SB0/n1296 ,
         \U1/aes_core/SB0/n1295 , \U1/aes_core/SB0/n1294 ,
         \U1/aes_core/SB0/n1293 , \U1/aes_core/SB0/n1292 ,
         \U1/aes_core/SB0/n1291 , \U1/aes_core/SB0/n1290 ,
         \U1/aes_core/SB0/n1289 , \U1/aes_core/SB0/n1288 ,
         \U1/aes_core/SB0/n1287 , \U1/aes_core/SB0/n1286 ,
         \U1/aes_core/SB0/n1285 , \U1/aes_core/SB0/n1284 ,
         \U1/aes_core/SB0/n1283 , \U1/aes_core/SB0/n1282 ,
         \U1/aes_core/SB0/n1281 , \U1/aes_core/SB0/n1280 ,
         \U1/aes_core/SB0/n1279 , \U1/aes_core/SB0/n1278 ,
         \U1/aes_core/SB0/n1277 , \U1/aes_core/SB0/n1276 ,
         \U1/aes_core/SB0/n1275 , \U1/aes_core/SB0/n1274 ,
         \U1/aes_core/SB0/n1273 , \U1/aes_core/SB0/n1272 ,
         \U1/aes_core/SB0/n1271 , \U1/aes_core/SB0/n1270 ,
         \U1/aes_core/SB0/n1269 , \U1/aes_core/SB0/n1268 ,
         \U1/aes_core/SB0/n1267 , \U1/aes_core/SB0/n1266 ,
         \U1/aes_core/SB0/n1265 , \U1/aes_core/SB0/n1264 ,
         \U1/aes_core/SB0/n1263 , \U1/aes_core/SB0/n1262 ,
         \U1/aes_core/SB0/n1261 , \U1/aes_core/SB0/n1260 ,
         \U1/aes_core/SB0/n1259 , \U1/aes_core/SB0/n1258 ,
         \U1/aes_core/SB0/n1257 , \U1/aes_core/SB0/n1256 ,
         \U1/aes_core/SB0/n1255 , \U1/aes_core/SB0/n1254 ,
         \U1/aes_core/SB0/n1253 , \U1/aes_core/SB0/n1252 ,
         \U1/aes_core/SB0/n1251 , \U1/aes_core/SB0/n1250 ,
         \U1/aes_core/SB0/n1249 , \U1/aes_core/SB0/n1248 ,
         \U1/aes_core/SB0/n1247 , \U1/aes_core/SB0/n1246 ,
         \U1/aes_core/SB0/n1245 , \U1/aes_core/SB0/n1244 ,
         \U1/aes_core/SB0/n1243 , \U1/aes_core/SB0/n1242 ,
         \U1/aes_core/SB0/n1241 , \U1/aes_core/SB0/n1240 ,
         \U1/aes_core/SB0/n1239 , \U1/aes_core/SB0/n1238 ,
         \U1/aes_core/SB0/n1237 , \U1/aes_core/SB0/n1236 ,
         \U1/aes_core/SB0/n1235 , \U1/aes_core/SB0/n1234 ,
         \U1/aes_core/SB0/n1233 , \U1/aes_core/SB0/n1232 ,
         \U1/aes_core/SB0/n1231 , \U1/aes_core/SB0/n1230 ,
         \U1/aes_core/SB0/n1229 , \U1/aes_core/SB0/n1228 ,
         \U1/aes_core/SB0/n1227 , \U1/aes_core/SB0/n1226 ,
         \U1/aes_core/SB0/n1225 , \U1/aes_core/SB0/n1224 ,
         \U1/aes_core/SB0/n1223 , \U1/aes_core/SB0/n1222 ,
         \U1/aes_core/SB0/n1221 , \U1/aes_core/SB0/n1220 ,
         \U1/aes_core/SB0/n1219 , \U1/aes_core/SB0/n1217 ,
         \U1/aes_core/SB0/n1216 , \U1/aes_core/SB0/n1215 ,
         \U1/aes_core/SB0/n1214 , \U1/aes_core/SB0/n1213 ,
         \U1/aes_core/SB0/n1212 , \U1/aes_core/SB0/n1211 ,
         \U1/aes_core/SB0/n1210 , \U1/aes_core/SB0/n1209 ,
         \U1/aes_core/SB0/n1208 , \U1/aes_core/SB0/n1207 ,
         \U1/aes_core/SB0/n1206 , \U1/aes_core/SB0/n1205 ,
         \U1/aes_core/SB0/n1204 , \U1/aes_core/SB0/n1202 ,
         \U1/aes_core/SB0/n1201 , \U1/aes_core/SB0/n1200 ,
         \U1/aes_core/SB0/n1199 , \U1/aes_core/SB0/n1198 ,
         \U1/aes_core/SB0/n1197 , \U1/aes_core/SB0/n1196 ,
         \U1/aes_core/SB0/n1195 , \U1/aes_core/SB0/n1194 ,
         \U1/aes_core/SB0/n1193 , \U1/aes_core/SB0/n1192 ,
         \U1/aes_core/SB0/n1191 , \U1/aes_core/SB0/n1190 ,
         \U1/aes_core/SB0/n1189 , \U1/aes_core/SB0/n1188 ,
         \U1/aes_core/SB0/n1187 , \U1/aes_core/SB0/n1186 ,
         \U1/aes_core/SB0/n1185 , \U1/aes_core/SB0/n1184 ,
         \U1/aes_core/SB0/n1183 , \U1/aes_core/SB0/n1182 ,
         \U1/aes_core/SB0/n1181 , \U1/aes_core/SB0/n1180 ,
         \U1/aes_core/SB0/n1179 , \U1/aes_core/SB0/n1178 ,
         \U1/aes_core/SB0/n1177 , \U1/aes_core/SB0/n1176 ,
         \U1/aes_core/SB0/n1175 , \U1/aes_core/SB0/n1174 ,
         \U1/aes_core/SB0/n1173 , \U1/aes_core/SB0/n1172 ,
         \U1/aes_core/SB0/n1171 , \U1/aes_core/SB0/n1170 ,
         \U1/aes_core/SB0/n1169 , \U1/aes_core/SB0/n1168 ,
         \U1/aes_core/SB0/n1167 , \U1/aes_core/SB0/n1166 ,
         \U1/aes_core/SB0/n1165 , \U1/aes_core/SB0/n1164 ,
         \U1/aes_core/SB0/n1163 , \U1/aes_core/SB0/n1162 ,
         \U1/aes_core/SB0/n1161 , \U1/aes_core/SB0/n1160 ,
         \U1/aes_core/SB0/n1159 , \U1/aes_core/SB0/n1157 ,
         \U1/aes_core/SB0/n1156 , \U1/aes_core/SB0/n1155 ,
         \U1/aes_core/SB0/n1154 , \U1/aes_core/SB0/n1153 ,
         \U1/aes_core/SB0/n1152 , \U1/aes_core/SB0/n1151 ,
         \U1/aes_core/SB0/n1150 , \U1/aes_core/SB0/n1149 ,
         \U1/aes_core/SB0/n1148 , \U1/aes_core/SB0/n1147 ,
         \U1/aes_core/SB0/n1146 , \U1/aes_core/SB0/n1145 ,
         \U1/aes_core/SB0/n1144 , \U1/aes_core/SB0/n1143 ,
         \U1/aes_core/SB0/n1142 , \U1/aes_core/SB0/n1141 ,
         \U1/aes_core/SB0/n1140 , \U1/aes_core/SB0/n1139 ,
         \U1/aes_core/SB0/n1138 , \U1/aes_core/SB0/n1137 ,
         \U1/aes_core/SB0/n1136 , \U1/aes_core/SB0/n1135 ,
         \U1/aes_core/SB0/n1134 , \U1/aes_core/SB0/n1133 ,
         \U1/aes_core/SB0/n1132 , \U1/aes_core/SB0/n1131 ,
         \U1/aes_core/SB0/n1130 , \U1/aes_core/SB0/n1129 ,
         \U1/aes_core/SB0/n1128 , \U1/aes_core/SB0/n1127 ,
         \U1/aes_core/SB0/n1126 , \U1/aes_core/SB0/n1125 ,
         \U1/aes_core/SB0/n1124 , \U1/aes_core/SB0/n1123 ,
         \U1/aes_core/SB0/n1122 , \U1/aes_core/SB0/n1121 ,
         \U1/aes_core/SB0/n1120 , \U1/aes_core/SB0/n1119 ,
         \U1/aes_core/SB0/n1118 , \U1/aes_core/SB0/n1117 ,
         \U1/aes_core/SB0/n1116 , \U1/aes_core/SB0/n1115 ,
         \U1/aes_core/SB0/n1114 , \U1/aes_core/SB0/n1113 ,
         \U1/aes_core/SB0/n1112 , \U1/aes_core/SB0/n1111 ,
         \U1/aes_core/SB0/n1110 , \U1/aes_core/SB0/n1109 ,
         \U1/aes_core/SB0/n1108 , \U1/aes_core/SB0/n1107 ,
         \U1/aes_core/SB0/n1106 , \U1/aes_core/SB0/n1105 ,
         \U1/aes_core/SB0/n1104 , \U1/aes_core/SB0/n1103 ,
         \U1/aes_core/SB0/n1102 , \U1/aes_core/SB0/n1101 ,
         \U1/aes_core/SB0/n1100 , \U1/aes_core/SB0/n1099 ,
         \U1/aes_core/SB0/n1098 , \U1/aes_core/SB0/n1097 ,
         \U1/aes_core/SB0/n1096 , \U1/aes_core/SB0/n1095 ,
         \U1/aes_core/SB0/n1094 , \U1/aes_core/SB0/n1093 ,
         \U1/aes_core/SB0/n1092 , \U1/aes_core/SB0/n1091 ,
         \U1/aes_core/SB0/n1090 , \U1/aes_core/SB0/n1089 ,
         \U1/aes_core/SB0/n1088 , \U1/aes_core/SB0/n1087 ,
         \U1/aes_core/SB0/n1086 , \U1/aes_core/SB0/n1085 ,
         \U1/aes_core/SB0/n1084 , \U1/aes_core/SB0/n1083 ,
         \U1/aes_core/SB0/n1082 , \U1/aes_core/SB0/n1081 ,
         \U1/aes_core/SB0/n1080 , \U1/aes_core/SB0/n1079 ,
         \U1/aes_core/SB0/n1078 , \U1/aes_core/SB0/n1077 ,
         \U1/aes_core/SB0/n1076 , \U1/aes_core/SB0/n1075 ,
         \U1/aes_core/SB0/n1074 , \U1/aes_core/SB0/n1073 ,
         \U1/aes_core/SB0/n1072 , \U1/aes_core/SB0/n1071 ,
         \U1/aes_core/SB0/n1070 , \U1/aes_core/SB0/n1069 ,
         \U1/aes_core/SB0/n1068 , \U1/aes_core/SB0/n1067 ,
         \U1/aes_core/SB0/n1066 , \U1/aes_core/SB0/n1065 ,
         \U1/aes_core/SB0/n1064 , \U1/aes_core/SB0/n1063 ,
         \U1/aes_core/SB0/n1062 , \U1/aes_core/SB0/n1061 ,
         \U1/aes_core/SB0/n1060 , \U1/aes_core/SB0/n1059 ,
         \U1/aes_core/SB0/n1058 , \U1/aes_core/SB0/n1057 ,
         \U1/aes_core/SB0/n1056 , \U1/aes_core/SB0/n1055 ,
         \U1/aes_core/SB0/n1054 , \U1/aes_core/SB0/n1053 ,
         \U1/aes_core/SB0/n1052 , \U1/aes_core/SB0/n1051 ,
         \U1/aes_core/SB0/n1050 , \U1/aes_core/SB0/n1049 ,
         \U1/aes_core/SB0/n1048 , \U1/aes_core/SB0/n1047 ,
         \U1/aes_core/SB0/n1046 , \U1/aes_core/SB0/n1045 ,
         \U1/aes_core/SB0/n1044 , \U1/aes_core/SB0/n1043 ,
         \U1/aes_core/SB0/n1042 , \U1/aes_core/SB0/n1041 ,
         \U1/aes_core/SB0/n1040 , \U1/aes_core/SB0/n1039 ,
         \U1/aes_core/SB0/n1038 , \U1/aes_core/SB0/n1037 ,
         \U1/aes_core/SB0/n1036 , \U1/aes_core/SB0/n1035 ,
         \U1/aes_core/SB0/n1034 , \U1/aes_core/SB0/n1033 ,
         \U1/aes_core/SB0/n1032 , \U1/aes_core/SB0/n1031 ,
         \U1/aes_core/SB0/n1029 , \U1/aes_core/SB0/n1028 ,
         \U1/aes_core/SB0/n1027 , \U1/aes_core/SB0/n1026 ,
         \U1/aes_core/SB0/n1025 , \U1/aes_core/SB0/n1024 ,
         \U1/aes_core/SB0/n1023 , \U1/aes_core/SB0/n1022 ,
         \U1/aes_core/SB0/n1021 , \U1/aes_core/SB0/n1020 ,
         \U1/aes_core/SB0/n1019 , \U1/aes_core/SB0/n1018 ,
         \U1/aes_core/SB0/n1017 , \U1/aes_core/SB0/n1016 ,
         \U1/aes_core/SB0/n1015 , \U1/aes_core/SB0/n1014 ,
         \U1/aes_core/SB0/n1013 , \U1/aes_core/SB0/n1012 ,
         \U1/aes_core/SB0/n1011 , \U1/aes_core/SB0/n1010 ,
         \U1/aes_core/SB0/n1009 , \U1/aes_core/SB0/n1008 ,
         \U1/aes_core/SB0/n1007 , \U1/aes_core/SB0/n1006 ,
         \U1/aes_core/SB0/n1005 , \U1/aes_core/SB0/n1004 ,
         \U1/aes_core/SB0/n1003 , \U1/aes_core/SB0/n1002 ,
         \U1/aes_core/SB0/n1001 , \U1/aes_core/SB0/n1000 ,
         \U1/aes_core/SB0/n999 , \U1/aes_core/SB0/n998 ,
         \U1/aes_core/SB0/n997 , \U1/aes_core/SB0/n996 ,
         \U1/aes_core/SB0/n995 , \U1/aes_core/SB0/n994 ,
         \U1/aes_core/SB0/n993 , \U1/aes_core/SB0/n992 ,
         \U1/aes_core/SB0/n991 , \U1/aes_core/SB0/n990 ,
         \U1/aes_core/SB0/n989 , \U1/aes_core/SB0/n988 ,
         \U1/aes_core/SB0/n987 , \U1/aes_core/SB0/n986 ,
         \U1/aes_core/SB0/n985 , \U1/aes_core/SB0/n984 ,
         \U1/aes_core/SB0/n983 , \U1/aes_core/SB0/n982 ,
         \U1/aes_core/SB0/n981 , \U1/aes_core/SB0/n980 ,
         \U1/aes_core/SB0/n979 , \U1/aes_core/SB0/n978 ,
         \U1/aes_core/SB0/n977 , \U1/aes_core/SB0/n976 ,
         \U1/aes_core/SB0/n975 , \U1/aes_core/SB0/n974 ,
         \U1/aes_core/SB0/n973 , \U1/aes_core/SB0/n972 ,
         \U1/aes_core/SB0/n971 , \U1/aes_core/SB0/n970 ,
         \U1/aes_core/SB0/n969 , \U1/aes_core/SB0/n968 ,
         \U1/aes_core/SB0/n967 , \U1/aes_core/SB0/n966 ,
         \U1/aes_core/SB0/n965 , \U1/aes_core/SB0/n964 ,
         \U1/aes_core/SB0/n963 , \U1/aes_core/SB0/n962 ,
         \U1/aes_core/SB0/n961 , \U1/aes_core/SB0/n960 ,
         \U1/aes_core/SB0/n959 , \U1/aes_core/SB0/n958 ,
         \U1/aes_core/SB0/n957 , \U1/aes_core/SB0/n956 ,
         \U1/aes_core/SB0/n955 , \U1/aes_core/SB0/n954 ,
         \U1/aes_core/SB0/n953 , \U1/aes_core/SB0/n952 ,
         \U1/aes_core/SB0/n951 , \U1/aes_core/SB0/n950 ,
         \U1/aes_core/SB0/n949 , \U1/aes_core/SB0/n948 ,
         \U1/aes_core/SB0/n947 , \U1/aes_core/SB0/n946 ,
         \U1/aes_core/SB0/n945 , \U1/aes_core/SB0/n944 ,
         \U1/aes_core/SB0/n943 , \U1/aes_core/SB0/n942 ,
         \U1/aes_core/SB0/n941 , \U1/aes_core/SB0/n940 ,
         \U1/aes_core/SB0/n939 , \U1/aes_core/SB0/n938 ,
         \U1/aes_core/SB0/n937 , \U1/aes_core/SB0/n936 ,
         \U1/aes_core/SB0/n935 , \U1/aes_core/SB0/n934 ,
         \U1/aes_core/SB0/n933 , \U1/aes_core/SB0/n932 ,
         \U1/aes_core/SB0/n931 , \U1/aes_core/SB0/n930 ,
         \U1/aes_core/SB0/n929 , \U1/aes_core/SB0/n928 ,
         \U1/aes_core/SB0/n927 , \U1/aes_core/SB0/n926 ,
         \U1/aes_core/SB0/n925 , \U1/aes_core/SB0/n924 ,
         \U1/aes_core/SB0/n923 , \U1/aes_core/SB0/n922 ,
         \U1/aes_core/SB0/n921 , \U1/aes_core/SB0/n920 ,
         \U1/aes_core/SB0/n919 , \U1/aes_core/SB0/n918 ,
         \U1/aes_core/SB0/n917 , \U1/aes_core/SB0/n916 ,
         \U1/aes_core/SB0/n915 , \U1/aes_core/SB0/n914 ,
         \U1/aes_core/SB0/n913 , \U1/aes_core/SB0/n912 ,
         \U1/aes_core/SB0/n911 , \U1/aes_core/SB0/n910 ,
         \U1/aes_core/SB0/n909 , \U1/aes_core/SB0/n908 ,
         \U1/aes_core/SB0/n907 , \U1/aes_core/SB0/n906 ,
         \U1/aes_core/SB0/n905 , \U1/aes_core/SB0/n904 ,
         \U1/aes_core/SB0/n903 , \U1/aes_core/SB0/n902 ,
         \U1/aes_core/SB0/n901 , \U1/aes_core/SB0/n900 ,
         \U1/aes_core/SB0/n899 , \U1/aes_core/SB0/n898 ,
         \U1/aes_core/SB0/n897 , \U1/aes_core/SB0/n896 ,
         \U1/aes_core/SB0/n895 , \U1/aes_core/SB0/n894 ,
         \U1/aes_core/SB0/n893 , \U1/aes_core/SB0/n892 ,
         \U1/aes_core/SB0/n891 , \U1/aes_core/SB0/n890 ,
         \U1/aes_core/SB0/n889 , \U1/aes_core/SB0/n888 ,
         \U1/aes_core/SB0/n887 , \U1/aes_core/SB0/n886 ,
         \U1/aes_core/SB0/n885 , \U1/aes_core/SB0/n884 ,
         \U1/aes_core/SB0/n883 , \U1/aes_core/SB0/n882 ,
         \U1/aes_core/SB0/n881 , \U1/aes_core/SB0/n880 ,
         \U1/aes_core/SB0/n879 , \U1/aes_core/SB0/n878 ,
         \U1/aes_core/SB0/n877 , \U1/aes_core/SB0/n876 ,
         \U1/aes_core/SB0/n875 , \U1/aes_core/SB0/n874 ,
         \U1/aes_core/SB0/n873 , \U1/aes_core/SB0/n872 ,
         \U1/aes_core/SB0/n871 , \U1/aes_core/SB0/n870 ,
         \U1/aes_core/SB0/n869 , \U1/aes_core/SB0/n868 ,
         \U1/aes_core/SB0/n867 , \U1/aes_core/SB0/n866 ,
         \U1/aes_core/SB0/n865 , \U1/aes_core/SB0/n864 ,
         \U1/aes_core/SB0/n863 , \U1/aes_core/SB0/n862 ,
         \U1/aes_core/SB0/n861 , \U1/aes_core/SB0/n860 ,
         \U1/aes_core/SB0/n859 , \U1/aes_core/SB0/n858 ,
         \U1/aes_core/SB0/n857 , \U1/aes_core/SB0/n856 ,
         \U1/aes_core/SB0/n855 , \U1/aes_core/SB0/n854 ,
         \U1/aes_core/SB0/n853 , \U1/aes_core/SB0/n852 ,
         \U1/aes_core/SB0/n851 , \U1/aes_core/SB0/n850 ,
         \U1/aes_core/SB0/n849 , \U1/aes_core/SB0/n848 ,
         \U1/aes_core/SB0/n847 , \U1/aes_core/SB0/n846 ,
         \U1/aes_core/SB0/n845 , \U1/aes_core/SB0/n844 ,
         \U1/aes_core/SB0/n843 , \U1/aes_core/SB0/n842 ,
         \U1/aes_core/SB0/n841 , \U1/aes_core/SB0/n840 ,
         \U1/aes_core/SB0/n839 , \U1/aes_core/SB0/n838 ,
         \U1/aes_core/SB0/n837 , \U1/aes_core/SB0/n836 ,
         \U1/aes_core/SB0/n835 , \U1/aes_core/SB0/n834 ,
         \U1/aes_core/SB0/n833 , \U1/aes_core/SB0/n832 ,
         \U1/aes_core/SB0/n831 , \U1/aes_core/SB0/n830 ,
         \U1/aes_core/SB0/n829 , \U1/aes_core/SB0/n828 ,
         \U1/aes_core/SB0/n827 , \U1/aes_core/SB0/n826 ,
         \U1/aes_core/SB0/n825 , \U1/aes_core/SB0/n824 ,
         \U1/aes_core/SB0/n823 , \U1/aes_core/SB0/n822 ,
         \U1/aes_core/SB0/n821 , \U1/aes_core/SB0/n820 ,
         \U1/aes_core/SB0/n819 , \U1/aes_core/SB0/n818 ,
         \U1/aes_core/SB0/n817 , \U1/aes_core/SB0/n816 ,
         \U1/aes_core/SB0/n815 , \U1/aes_core/SB0/n814 ,
         \U1/aes_core/SB0/n813 , \U1/aes_core/SB0/n812 ,
         \U1/aes_core/SB0/n811 , \U1/aes_core/SB0/n810 ,
         \U1/aes_core/SB0/n809 , \U1/aes_core/SB0/n808 ,
         \U1/aes_core/SB0/n807 , \U1/aes_core/SB0/n806 ,
         \U1/aes_core/SB0/n805 , \U1/aes_core/SB0/n804 ,
         \U1/aes_core/SB0/n803 , \U1/aes_core/SB0/n802 ,
         \U1/aes_core/SB0/n801 , \U1/aes_core/SB0/n800 ,
         \U1/aes_core/SB0/n799 , \U1/aes_core/SB0/n798 ,
         \U1/aes_core/SB0/n797 , \U1/aes_core/SB0/n796 ,
         \U1/aes_core/SB0/n795 , \U1/aes_core/SB0/n794 ,
         \U1/aes_core/SB0/n793 , \U1/aes_core/SB0/n792 ,
         \U1/aes_core/SB0/n791 , \U1/aes_core/SB0/n790 ,
         \U1/aes_core/SB0/n789 , \U1/aes_core/SB0/n788 ,
         \U1/aes_core/SB0/n787 , \U1/aes_core/SB0/n786 ,
         \U1/aes_core/SB0/n785 , \U1/aes_core/SB0/n784 ,
         \U1/aes_core/SB0/n783 , \U1/aes_core/SB0/n782 ,
         \U1/aes_core/SB0/n781 , \U1/aes_core/SB0/n780 ,
         \U1/aes_core/SB0/n779 , \U1/aes_core/SB0/n778 ,
         \U1/aes_core/SB0/n777 , \U1/aes_core/SB0/n776 ,
         \U1/aes_core/SB0/n775 , \U1/aes_core/SB0/n774 ,
         \U1/aes_core/SB0/n773 , \U1/aes_core/SB0/n772 ,
         \U1/aes_core/SB0/n771 , \U1/aes_core/SB0/n770 ,
         \U1/aes_core/SB0/n769 , \U1/aes_core/SB0/n768 ,
         \U1/aes_core/SB0/n766 , \U1/aes_core/SB0/n765 ,
         \U1/aes_core/SB0/n764 , \U1/aes_core/SB0/n763 ,
         \U1/aes_core/SB0/n762 , \U1/aes_core/SB0/n761 ,
         \U1/aes_core/SB0/n760 , \U1/aes_core/SB0/n759 ,
         \U1/aes_core/SB0/n758 , \U1/aes_core/SB0/n757 ,
         \U1/aes_core/SB0/n756 , \U1/aes_core/SB0/n755 ,
         \U1/aes_core/SB0/n754 , \U1/aes_core/SB0/n753 ,
         \U1/aes_core/SB0/n751 , \U1/aes_core/SB0/n750 ,
         \U1/aes_core/SB0/n749 , \U1/aes_core/SB0/n748 ,
         \U1/aes_core/SB0/n747 , \U1/aes_core/SB0/n746 ,
         \U1/aes_core/SB0/n745 , \U1/aes_core/SB0/n744 ,
         \U1/aes_core/SB0/n743 , \U1/aes_core/SB0/n742 ,
         \U1/aes_core/SB0/n741 , \U1/aes_core/SB0/n740 ,
         \U1/aes_core/SB0/n739 , \U1/aes_core/SB0/n738 ,
         \U1/aes_core/SB0/n737 , \U1/aes_core/SB0/n736 ,
         \U1/aes_core/SB0/n735 , \U1/aes_core/SB0/n734 ,
         \U1/aes_core/SB0/n733 , \U1/aes_core/SB0/n732 ,
         \U1/aes_core/SB0/n731 , \U1/aes_core/SB0/n730 ,
         \U1/aes_core/SB0/n729 , \U1/aes_core/SB0/n728 ,
         \U1/aes_core/SB0/n727 , \U1/aes_core/SB0/n726 ,
         \U1/aes_core/SB0/n725 , \U1/aes_core/SB0/n724 ,
         \U1/aes_core/SB0/n723 , \U1/aes_core/SB0/n722 ,
         \U1/aes_core/SB0/n721 , \U1/aes_core/SB0/n720 ,
         \U1/aes_core/SB0/n719 , \U1/aes_core/SB0/n718 ,
         \U1/aes_core/SB0/n717 , \U1/aes_core/SB0/n716 ,
         \U1/aes_core/SB0/n715 , \U1/aes_core/SB0/n714 ,
         \U1/aes_core/SB0/n713 , \U1/aes_core/SB0/n712 ,
         \U1/aes_core/SB0/n711 , \U1/aes_core/SB0/n710 ,
         \U1/aes_core/SB0/n709 , \U1/aes_core/SB0/n708 ,
         \U1/aes_core/SB0/n706 , \U1/aes_core/SB0/n705 ,
         \U1/aes_core/SB0/n704 , \U1/aes_core/SB0/n703 ,
         \U1/aes_core/SB0/n702 , \U1/aes_core/SB0/n701 ,
         \U1/aes_core/SB0/n700 , \U1/aes_core/SB0/n699 ,
         \U1/aes_core/SB0/n698 , \U1/aes_core/SB0/n697 ,
         \U1/aes_core/SB0/n696 , \U1/aes_core/SB0/n695 ,
         \U1/aes_core/SB0/n694 , \U1/aes_core/SB0/n693 ,
         \U1/aes_core/SB0/n692 , \U1/aes_core/SB0/n691 ,
         \U1/aes_core/SB0/n690 , \U1/aes_core/SB0/n689 ,
         \U1/aes_core/SB0/n688 , \U1/aes_core/SB0/n687 ,
         \U1/aes_core/SB0/n686 , \U1/aes_core/SB0/n685 ,
         \U1/aes_core/SB0/n684 , \U1/aes_core/SB0/n683 ,
         \U1/aes_core/SB0/n682 , \U1/aes_core/SB0/n681 ,
         \U1/aes_core/SB0/n680 , \U1/aes_core/SB0/n679 ,
         \U1/aes_core/SB0/n678 , \U1/aes_core/SB0/n677 ,
         \U1/aes_core/SB0/n676 , \U1/aes_core/SB0/n675 ,
         \U1/aes_core/SB0/n674 , \U1/aes_core/SB0/n673 ,
         \U1/aes_core/SB0/n672 , \U1/aes_core/SB0/n671 ,
         \U1/aes_core/SB0/n670 , \U1/aes_core/SB0/n669 ,
         \U1/aes_core/SB0/n668 , \U1/aes_core/SB0/n667 ,
         \U1/aes_core/SB0/n666 , \U1/aes_core/SB0/n665 ,
         \U1/aes_core/SB0/n664 , \U1/aes_core/SB0/n663 ,
         \U1/aes_core/SB0/n662 , \U1/aes_core/SB0/n661 ,
         \U1/aes_core/SB0/n660 , \U1/aes_core/SB0/n659 ,
         \U1/aes_core/SB0/n658 , \U1/aes_core/SB0/n657 ,
         \U1/aes_core/SB0/n656 , \U1/aes_core/SB0/n655 ,
         \U1/aes_core/SB0/n654 , \U1/aes_core/SB0/n653 ,
         \U1/aes_core/SB0/n652 , \U1/aes_core/SB0/n651 ,
         \U1/aes_core/SB0/n650 , \U1/aes_core/SB0/n649 ,
         \U1/aes_core/SB0/n648 , \U1/aes_core/SB0/n647 ,
         \U1/aes_core/SB0/n646 , \U1/aes_core/SB0/n645 ,
         \U1/aes_core/SB0/n644 , \U1/aes_core/SB0/n643 ,
         \U1/aes_core/SB0/n642 , \U1/aes_core/SB0/n641 ,
         \U1/aes_core/SB0/n640 , \U1/aes_core/SB0/n639 ,
         \U1/aes_core/SB0/n638 , \U1/aes_core/SB0/n637 ,
         \U1/aes_core/SB0/n636 , \U1/aes_core/SB0/n635 ,
         \U1/aes_core/SB0/n634 , \U1/aes_core/SB0/n633 ,
         \U1/aes_core/SB0/n632 , \U1/aes_core/SB0/n631 ,
         \U1/aes_core/SB0/n630 , \U1/aes_core/SB0/n629 ,
         \U1/aes_core/SB0/n628 , \U1/aes_core/SB0/n627 ,
         \U1/aes_core/SB0/n626 , \U1/aes_core/SB0/n625 ,
         \U1/aes_core/SB0/n624 , \U1/aes_core/SB0/n623 ,
         \U1/aes_core/SB0/n622 , \U1/aes_core/SB0/n621 ,
         \U1/aes_core/SB0/n620 , \U1/aes_core/SB0/n619 ,
         \U1/aes_core/SB0/n618 , \U1/aes_core/SB0/n617 ,
         \U1/aes_core/SB0/n616 , \U1/aes_core/SB0/n615 ,
         \U1/aes_core/SB0/n614 , \U1/aes_core/SB0/n613 ,
         \U1/aes_core/SB0/n612 , \U1/aes_core/SB0/n611 ,
         \U1/aes_core/SB0/n610 , \U1/aes_core/SB0/n609 ,
         \U1/aes_core/SB0/n608 , \U1/aes_core/SB0/n607 ,
         \U1/aes_core/SB0/n606 , \U1/aes_core/SB0/n605 ,
         \U1/aes_core/SB0/n604 , \U1/aes_core/SB0/n603 ,
         \U1/aes_core/SB0/n602 , \U1/aes_core/SB0/n601 ,
         \U1/aes_core/SB0/n600 , \U1/aes_core/SB0/n599 ,
         \U1/aes_core/SB0/n598 , \U1/aes_core/SB0/n597 ,
         \U1/aes_core/SB0/n596 , \U1/aes_core/SB0/n595 ,
         \U1/aes_core/SB0/n594 , \U1/aes_core/SB0/n593 ,
         \U1/aes_core/SB0/n592 , \U1/aes_core/SB0/n591 ,
         \U1/aes_core/SB0/n590 , \U1/aes_core/SB0/n589 ,
         \U1/aes_core/SB0/n588 , \U1/aes_core/SB0/n587 ,
         \U1/aes_core/SB0/n586 , \U1/aes_core/SB0/n585 ,
         \U1/aes_core/SB0/n584 , \U1/aes_core/SB0/n583 ,
         \U1/aes_core/SB0/n582 , \U1/aes_core/SB0/n581 ,
         \U1/aes_core/SB0/n580 , \U1/aes_core/SB0/n579 ,
         \U1/aes_core/SB0/n578 , \U1/aes_core/SB0/n577 ,
         \U1/aes_core/SB0/n576 , \U1/aes_core/SB0/n575 ,
         \U1/aes_core/SB0/n574 , \U1/aes_core/SB0/n573 ,
         \U1/aes_core/SB0/n572 , \U1/aes_core/SB0/n571 ,
         \U1/aes_core/SB0/n570 , \U1/aes_core/SB0/n569 ,
         \U1/aes_core/SB0/n568 , \U1/aes_core/SB0/n567 ,
         \U1/aes_core/SB0/n566 , \U1/aes_core/SB0/n565 ,
         \U1/aes_core/SB0/n564 , \U1/aes_core/SB0/n563 ,
         \U1/aes_core/SB0/n562 , \U1/aes_core/SB0/n561 ,
         \U1/aes_core/SB0/n560 , \U1/aes_core/SB0/n559 ,
         \U1/aes_core/SB0/n558 , \U1/aes_core/SB0/n557 ,
         \U1/aes_core/SB0/n556 , \U1/aes_core/SB0/n555 ,
         \U1/aes_core/SB0/n554 , \U1/aes_core/SB0/n553 ,
         \U1/aes_core/SB0/n552 , \U1/aes_core/SB0/n551 ,
         \U1/aes_core/SB0/n550 , \U1/aes_core/SB0/n549 ,
         \U1/aes_core/SB0/n548 , \U1/aes_core/SB0/n547 ,
         \U1/aes_core/SB0/n546 , \U1/aes_core/SB0/n545 ,
         \U1/aes_core/SB0/n544 , \U1/aes_core/SB0/n543 ,
         \U1/aes_core/SB0/n542 , \U1/aes_core/SB0/n541 ,
         \U1/aes_core/SB0/n540 , \U1/aes_core/SB0/n539 ,
         \U1/aes_core/SB0/n538 , \U1/aes_core/SB0/n537 ,
         \U1/aes_core/SB0/n536 , \U1/aes_core/SB0/n535 ,
         \U1/aes_core/SB0/n534 , \U1/aes_core/SB0/n533 ,
         \U1/aes_core/SB0/n532 , \U1/aes_core/SB0/n531 ,
         \U1/aes_core/SB0/n530 , \U1/aes_core/SB0/n529 ,
         \U1/aes_core/SB0/n528 , \U1/aes_core/SB0/n527 ,
         \U1/aes_core/SB0/n526 , \U1/aes_core/SB0/n525 ,
         \U1/aes_core/SB0/n524 , \U1/aes_core/SB0/n523 ,
         \U1/aes_core/SB0/n522 , \U1/aes_core/SB0/n521 ,
         \U1/aes_core/SB0/n520 , \U1/aes_core/SB0/n519 ,
         \U1/aes_core/SB0/n518 , \U1/aes_core/SB0/n517 ,
         \U1/aes_core/SB0/n516 , \U1/aes_core/SB0/n515 ,
         \U1/aes_core/SB0/n514 , \U1/aes_core/SB0/n513 ,
         \U1/aes_core/SB0/n512 , \U1/aes_core/SB0/n511 ,
         \U1/aes_core/SB0/n510 , \U1/aes_core/SB0/n509 ,
         \U1/aes_core/SB0/n508 , \U1/aes_core/SB0/n507 ,
         \U1/aes_core/SB0/n506 , \U1/aes_core/SB0/n505 ,
         \U1/aes_core/SB0/n504 , \U1/aes_core/SB0/n503 ,
         \U1/aes_core/SB0/n502 , \U1/aes_core/SB0/n501 ,
         \U1/aes_core/SB0/n500 , \U1/aes_core/SB0/n499 ,
         \U1/aes_core/SB0/n498 , \U1/aes_core/SB0/n497 ,
         \U1/aes_core/SB0/n496 , \U1/aes_core/SB0/n495 ,
         \U1/aes_core/SB0/n494 , \U1/aes_core/SB0/n493 ,
         \U1/aes_core/SB0/n492 , \U1/aes_core/SB0/n491 ,
         \U1/aes_core/SB0/n490 , \U1/aes_core/SB0/n489 ,
         \U1/aes_core/SB0/n488 , \U1/aes_core/SB0/n487 ,
         \U1/aes_core/SB0/n486 , \U1/aes_core/SB0/n485 ,
         \U1/aes_core/SB0/n484 , \U1/aes_core/SB0/n483 ,
         \U1/aes_core/SB0/n482 , \U1/aes_core/SB0/n481 ,
         \U1/aes_core/SB0/n480 , \U1/aes_core/SB0/n479 ,
         \U1/aes_core/SB0/n478 , \U1/aes_core/SB0/n477 ,
         \U1/aes_core/SB0/n476 , \U1/aes_core/SB0/n475 ,
         \U1/aes_core/SB0/n474 , \U1/aes_core/SB0/n473 ,
         \U1/aes_core/SB0/n472 , \U1/aes_core/SB0/n471 ,
         \U1/aes_core/SB0/n470 , \U1/aes_core/SB0/n469 ,
         \U1/aes_core/SB0/n468 , \U1/aes_core/SB0/n467 ,
         \U1/aes_core/SB0/n466 , \U1/aes_core/SB0/n465 ,
         \U1/aes_core/SB0/n464 , \U1/aes_core/SB0/n463 ,
         \U1/aes_core/SB0/n462 , \U1/aes_core/SB0/n461 ,
         \U1/aes_core/SB0/n460 , \U1/aes_core/SB0/n459 ,
         \U1/aes_core/SB0/n458 , \U1/aes_core/SB0/n457 ,
         \U1/aes_core/SB0/n456 , \U1/aes_core/SB0/n455 ,
         \U1/aes_core/SB0/n454 , \U1/aes_core/SB0/n453 ,
         \U1/aes_core/SB0/n452 , \U1/aes_core/SB0/n451 ,
         \U1/aes_core/SB0/n450 , \U1/aes_core/SB0/n449 ,
         \U1/aes_core/SB0/n448 , \U1/aes_core/SB0/n447 ,
         \U1/aes_core/SB0/n446 , \U1/aes_core/SB0/n445 ,
         \U1/aes_core/SB0/n444 , \U1/aes_core/SB0/n443 ,
         \U1/aes_core/SB0/n442 , \U1/aes_core/SB0/n441 ,
         \U1/aes_core/SB0/n440 , \U1/aes_core/SB0/n439 ,
         \U1/aes_core/SB0/n438 , \U1/aes_core/SB0/n437 ,
         \U1/aes_core/SB0/n436 , \U1/aes_core/SB0/n435 ,
         \U1/aes_core/SB0/n434 , \U1/aes_core/SB0/n433 ,
         \U1/aes_core/SB0/n432 , \U1/aes_core/SB0/n431 ,
         \U1/aes_core/SB0/n430 , \U1/aes_core/SB0/n429 ,
         \U1/aes_core/SB0/n428 , \U1/aes_core/SB0/n427 ,
         \U1/aes_core/SB0/n426 , \U1/aes_core/SB0/n425 ,
         \U1/aes_core/SB0/n424 , \U1/aes_core/SB0/n423 ,
         \U1/aes_core/SB0/n422 , \U1/aes_core/SB0/n421 ,
         \U1/aes_core/SB0/n420 , \U1/aes_core/SB0/n419 ,
         \U1/aes_core/SB0/n418 , \U1/aes_core/SB0/n417 ,
         \U1/aes_core/SB0/n416 , \U1/aes_core/SB0/n415 ,
         \U1/aes_core/SB0/n414 , \U1/aes_core/SB0/n413 ,
         \U1/aes_core/SB0/n412 , \U1/aes_core/SB0/n411 ,
         \U1/aes_core/SB0/n410 , \U1/aes_core/SB0/n409 ,
         \U1/aes_core/SB0/n408 , \U1/aes_core/SB0/n407 ,
         \U1/aes_core/SB0/n406 , \U1/aes_core/SB0/n405 ,
         \U1/aes_core/SB0/n404 , \U1/aes_core/SB0/n403 ,
         \U1/aes_core/SB0/n402 , \U1/aes_core/SB0/n401 ,
         \U1/aes_core/SB0/n400 , \U1/aes_core/SB0/n399 ,
         \U1/aes_core/SB0/n398 , \U1/aes_core/SB0/n397 ,
         \U1/aes_core/SB0/n396 , \U1/aes_core/SB0/n395 ,
         \U1/aes_core/SB0/n394 , \U1/aes_core/SB0/n393 ,
         \U1/aes_core/SB0/n392 , \U1/aes_core/SB0/n391 ,
         \U1/aes_core/SB0/n390 , \U1/aes_core/SB0/n389 ,
         \U1/aes_core/SB0/n388 , \U1/aes_core/SB0/n387 ,
         \U1/aes_core/SB0/n386 , \U1/aes_core/SB0/n384 ,
         \U1/aes_core/SB0/n383 , \U1/aes_core/SB0/n382 ,
         \U1/aes_core/SB0/n381 , \U1/aes_core/SB0/n380 ,
         \U1/aes_core/SB0/n379 , \U1/aes_core/SB0/n378 ,
         \U1/aes_core/SB0/n377 , \U1/aes_core/SB0/n376 ,
         \U1/aes_core/SB0/n375 , \U1/aes_core/SB0/n374 ,
         \U1/aes_core/SB0/n373 , \U1/aes_core/SB0/n372 ,
         \U1/aes_core/SB0/n371 , \U1/aes_core/SB0/n370 ,
         \U1/aes_core/SB0/n369 , \U1/aes_core/SB0/n368 ,
         \U1/aes_core/SB0/n367 , \U1/aes_core/SB0/n366 ,
         \U1/aes_core/SB0/n365 , \U1/aes_core/SB0/n364 ,
         \U1/aes_core/SB0/n363 , \U1/aes_core/SB0/n362 ,
         \U1/aes_core/SB0/n361 , \U1/aes_core/SB0/n360 ,
         \U1/aes_core/SB0/n359 , \U1/aes_core/SB0/n358 ,
         \U1/aes_core/SB0/n357 , \U1/aes_core/SB0/n356 ,
         \U1/aes_core/SB0/n355 , \U1/aes_core/SB0/n354 ,
         \U1/aes_core/SB0/n353 , \U1/aes_core/SB0/n352 ,
         \U1/aes_core/SB0/n351 , \U1/aes_core/SB0/n350 ,
         \U1/aes_core/SB0/n349 , \U1/aes_core/SB0/n348 ,
         \U1/aes_core/SB0/n347 , \U1/aes_core/SB0/n346 ,
         \U1/aes_core/SB0/n345 , \U1/aes_core/SB0/n344 ,
         \U1/aes_core/SB0/n343 , \U1/aes_core/SB0/n342 ,
         \U1/aes_core/SB0/n341 , \U1/aes_core/SB0/n340 ,
         \U1/aes_core/SB0/n339 , \U1/aes_core/SB0/n338 ,
         \U1/aes_core/SB0/n337 , \U1/aes_core/SB0/n336 ,
         \U1/aes_core/SB0/n335 , \U1/aes_core/SB0/n334 ,
         \U1/aes_core/SB0/n333 , \U1/aes_core/SB0/n332 ,
         \U1/aes_core/SB0/n331 , \U1/aes_core/SB0/n330 ,
         \U1/aes_core/SB0/n329 , \U1/aes_core/SB0/n328 ,
         \U1/aes_core/SB0/n327 , \U1/aes_core/SB0/n326 ,
         \U1/aes_core/SB0/n325 , \U1/aes_core/SB0/n324 ,
         \U1/aes_core/SB0/n323 , \U1/aes_core/SB0/n322 ,
         \U1/aes_core/SB0/n321 , \U1/aes_core/SB0/n320 ,
         \U1/aes_core/SB0/n319 , \U1/aes_core/SB0/n318 ,
         \U1/aes_core/SB0/n317 , \U1/aes_core/SB0/n316 ,
         \U1/aes_core/SB0/n315 , \U1/aes_core/SB0/n314 ,
         \U1/aes_core/SB0/n313 , \U1/aes_core/SB0/n312 ,
         \U1/aes_core/SB0/n311 , \U1/aes_core/SB0/n310 ,
         \U1/aes_core/SB0/n309 , \U1/aes_core/SB0/n308 ,
         \U1/aes_core/SB0/n307 , \U1/aes_core/SB0/n306 ,
         \U1/aes_core/SB0/n305 , \U1/aes_core/SB0/n304 ,
         \U1/aes_core/SB0/n303 , \U1/aes_core/SB0/n302 ,
         \U1/aes_core/SB0/n301 , \U1/aes_core/SB0/n300 ,
         \U1/aes_core/SB0/n299 , \U1/aes_core/SB0/n298 ,
         \U1/aes_core/SB0/n297 , \U1/aes_core/SB0/n296 ,
         \U1/aes_core/SB0/n295 , \U1/aes_core/SB0/n294 ,
         \U1/aes_core/SB0/n293 , \U1/aes_core/SB0/n292 ,
         \U1/aes_core/SB0/n291 , \U1/aes_core/SB0/n290 ,
         \U1/aes_core/SB0/n289 , \U1/aes_core/SB0/n288 ,
         \U1/aes_core/SB0/n287 , \U1/aes_core/SB0/n286 ,
         \U1/aes_core/SB0/n285 , \U1/aes_core/SB0/n284 ,
         \U1/aes_core/SB0/n283 , \U1/aes_core/SB0/n282 ,
         \U1/aes_core/SB0/n281 , \U1/aes_core/SB0/n280 ,
         \U1/aes_core/SB0/n279 , \U1/aes_core/SB0/n278 ,
         \U1/aes_core/SB0/n277 , \U1/aes_core/SB0/n276 ,
         \U1/aes_core/SB0/n275 , \U1/aes_core/SB0/n274 ,
         \U1/aes_core/SB0/n273 , \U1/aes_core/SB0/n272 ,
         \U1/aes_core/SB0/n271 , \U1/aes_core/SB0/n270 ,
         \U1/aes_core/SB0/n269 , \U1/aes_core/SB0/n268 ,
         \U1/aes_core/SB0/n267 , \U1/aes_core/SB0/n266 ,
         \U1/aes_core/SB0/n265 , \U1/aes_core/SB0/n264 ,
         \U1/aes_core/SB0/n263 , \U1/aes_core/SB0/n262 ,
         \U1/aes_core/SB0/n261 , \U1/aes_core/SB0/n260 ,
         \U1/aes_core/SB0/n259 , \U1/aes_core/SB0/n258 ,
         \U1/aes_core/SB0/n257 , \U1/aes_core/SB0/n256 ,
         \U1/aes_core/SB0/n255 , \U1/aes_core/SB0/n254 ,
         \U1/aes_core/SB0/n253 , \U1/aes_core/SB0/n252 ,
         \U1/aes_core/SB0/n251 , \U1/aes_core/SB0/n250 ,
         \U1/aes_core/SB0/n249 , \U1/aes_core/SB0/n248 ,
         \U1/aes_core/SB0/n247 , \U1/aes_core/SB0/n246 ,
         \U1/aes_core/SB0/n245 , \U1/aes_core/SB0/n244 ,
         \U1/aes_core/SB0/n243 , \U1/aes_core/SB0/n242 ,
         \U1/aes_core/SB0/n241 , \U1/aes_core/SB0/n240 ,
         \U1/aes_core/SB0/n239 , \U1/aes_core/SB0/n238 ,
         \U1/aes_core/SB0/n237 , \U1/aes_core/SB0/n236 ,
         \U1/aes_core/SB0/n235 , \U1/aes_core/SB0/n234 ,
         \U1/aes_core/SB0/n233 , \U1/aes_core/SB0/n232 ,
         \U1/aes_core/SB0/n231 , \U1/aes_core/SB0/n230 ,
         \U1/aes_core/SB0/n229 , \U1/aes_core/SB0/n228 ,
         \U1/aes_core/SB0/n227 , \U1/aes_core/SB0/n226 ,
         \U1/aes_core/SB0/n225 , \U1/aes_core/SB0/n224 ,
         \U1/aes_core/SB0/n223 , \U1/aes_core/SB0/n222 ,
         \U1/aes_core/SB0/n221 , \U1/aes_core/SB0/n220 ,
         \U1/aes_core/SB0/n219 , \U1/aes_core/SB0/n218 ,
         \U1/aes_core/SB0/n217 , \U1/aes_core/SB0/n216 ,
         \U1/aes_core/SB0/n215 , \U1/aes_core/SB0/n214 ,
         \U1/aes_core/SB0/n213 , \U1/aes_core/SB0/n212 ,
         \U1/aes_core/SB0/n211 , \U1/aes_core/SB0/n210 ,
         \U1/aes_core/SB0/n209 , \U1/aes_core/SB0/n208 ,
         \U1/aes_core/SB0/n207 , \U1/aes_core/SB0/n206 ,
         \U1/aes_core/SB0/n205 , \U1/aes_core/SB0/n204 ,
         \U1/aes_core/SB0/n203 , \U1/aes_core/SB0/n202 ,
         \U1/aes_core/SB0/n201 , \U1/aes_core/SB0/n200 ,
         \U1/aes_core/SB0/n199 , \U1/aes_core/SB0/n198 ,
         \U1/aes_core/SB0/n197 , \U1/aes_core/SB0/n196 ,
         \U1/aes_core/SB0/n195 , \U1/aes_core/SB0/n194 ,
         \U1/aes_core/SB0/n193 , \U1/aes_core/SB0/n192 ,
         \U1/aes_core/SB0/n191 , \U1/aes_core/SB0/n190 ,
         \U1/aes_core/SB0/n189 , \U1/aes_core/SB0/n188 ,
         \U1/aes_core/SB0/n187 , \U1/aes_core/SB0/n186 ,
         \U1/aes_core/SB0/n185 , \U1/aes_core/SB0/n184 ,
         \U1/aes_core/SB0/n183 , \U1/aes_core/SB0/n182 ,
         \U1/aes_core/SB0/n181 , \U1/aes_core/SB0/n180 ,
         \U1/aes_core/SB0/n179 , \U1/aes_core/SB0/n178 ,
         \U1/aes_core/SB0/n177 , \U1/aes_core/SB0/n176 ,
         \U1/aes_core/SB0/n175 , \U1/aes_core/SB0/n174 ,
         \U1/aes_core/SB0/n173 , \U1/aes_core/SB0/n172 ,
         \U1/aes_core/SB0/n171 , \U1/aes_core/SB0/n170 ,
         \U1/aes_core/SB0/n169 , \U1/aes_core/SB0/n168 ,
         \U1/aes_core/SB0/n167 , \U1/aes_core/SB0/n166 ,
         \U1/aes_core/SB0/n165 , \U1/aes_core/SB0/n164 ,
         \U1/aes_core/SB0/n163 , \U1/aes_core/SB0/n162 ,
         \U1/aes_core/SB0/n161 , \U1/aes_core/SB0/n160 ,
         \U1/aes_core/SB0/n159 , \U1/aes_core/SB0/n158 ,
         \U1/aes_core/SB0/n157 , \U1/aes_core/SB0/n156 ,
         \U1/aes_core/SB0/n155 , \U1/aes_core/SB0/n154 ,
         \U1/aes_core/SB0/n153 , \U1/aes_core/SB0/n152 ,
         \U1/aes_core/SB0/n151 , \U1/aes_core/SB0/n150 ,
         \U1/aes_core/SB0/n149 , \U1/aes_core/SB0/n148 ,
         \U1/aes_core/SB0/n147 , \U1/aes_core/SB0/n146 ,
         \U1/aes_core/SB0/n145 , \U1/aes_core/SB0/n144 ,
         \U1/aes_core/SB0/n143 , \U1/aes_core/SB0/n142 ,
         \U1/aes_core/SB0/n141 , \U1/aes_core/SB0/n140 ,
         \U1/aes_core/SB0/n139 , \U1/aes_core/SB0/n138 ,
         \U1/aes_core/SB0/n137 , \U1/aes_core/SB0/n136 ,
         \U1/aes_core/SB0/n135 , \U1/aes_core/SB0/n134 ,
         \U1/aes_core/SB0/n133 , \U1/aes_core/SB0/n132 ,
         \U1/aes_core/SB0/n131 , \U1/aes_core/SB0/n130 ,
         \U1/aes_core/SB0/n129 , \U1/aes_core/SB0/n128 ,
         \U1/aes_core/SB0/n127 , \U1/aes_core/SB0/n126 ,
         \U1/aes_core/SB0/n125 , \U1/aes_core/SB0/n124 ,
         \U1/aes_core/SB0/n123 , \U1/aes_core/SB0/n122 ,
         \U1/aes_core/SB0/n121 , \U1/aes_core/SB0/n120 ,
         \U1/aes_core/SB0/n119 , \U1/aes_core/SB0/n118 ,
         \U1/aes_core/SB0/n117 , \U1/aes_core/SB0/n116 ,
         \U1/aes_core/SB0/n115 , \U1/aes_core/SB0/n114 ,
         \U1/aes_core/SB0/n113 , \U1/aes_core/SB0/n112 ,
         \U1/aes_core/SB0/n111 , \U1/aes_core/SB0/n110 ,
         \U1/aes_core/SB0/n109 , \U1/aes_core/SB0/n108 ,
         \U1/aes_core/SB0/n107 , \U1/aes_core/SB0/n106 ,
         \U1/aes_core/SB0/n105 , \U1/aes_core/SB0/n104 ,
         \U1/aes_core/SB0/n103 , \U1/aes_core/SB0/n102 ,
         \U1/aes_core/SB0/n101 , \U1/aes_core/SB0/n100 , \U1/aes_core/SB0/n99 ,
         \U1/aes_core/SB0/n98 , \U1/aes_core/SB0/n97 , \U1/aes_core/SB0/n96 ,
         \U1/aes_core/SB0/n95 , \U1/aes_core/SB0/n94 , \U1/aes_core/SB0/n93 ,
         \U1/aes_core/SB0/n92 , \U1/aes_core/SB0/n91 , \U1/aes_core/SB0/n90 ,
         \U1/aes_core/SB0/n89 , \U1/aes_core/SB0/n88 , \U1/aes_core/SB0/n87 ,
         \U1/aes_core/SB0/n86 , \U1/aes_core/SB0/n85 , \U1/aes_core/SB0/n84 ,
         \U1/aes_core/SB0/n83 , \U1/aes_core/SB0/n82 , \U1/aes_core/SB0/n81 ,
         \U1/aes_core/SB0/n80 , \U1/aes_core/SB0/n79 , \U1/aes_core/SB0/n78 ,
         \U1/aes_core/SB0/n77 , \U1/aes_core/SB0/n76 , \U1/aes_core/SB0/n75 ,
         \U1/aes_core/SB0/n74 , \U1/aes_core/SB0/n73 , \U1/aes_core/SB0/n72 ,
         \U1/aes_core/SB0/n71 , \U1/aes_core/SB0/n70 , \U1/aes_core/SB0/n69 ,
         \U1/aes_core/SB0/n68 , \U1/aes_core/SB0/n67 , \U1/aes_core/SB0/n66 ,
         \U1/aes_core/SB0/n65 , \U1/aes_core/SB0/n64 , \U1/aes_core/SB0/n63 ,
         \U1/aes_core/SB0/n62 , \U1/aes_core/SB0/n61 , \U1/aes_core/SB0/n60 ,
         \U1/aes_core/SB0/n59 , \U1/aes_core/SB0/n58 , \U1/aes_core/SB0/n57 ,
         \U1/aes_core/SB0/n56 , \U1/aes_core/SB0/n55 , \U1/aes_core/SB0/n54 ,
         \U1/aes_core/SB0/n53 , \U1/aes_core/SB0/n52 , \U1/aes_core/SB0/n51 ,
         \U1/aes_core/SB0/n50 , \U1/aes_core/SB0/n49 , \U1/aes_core/SB0/n48 ,
         \U1/aes_core/SB0/n47 , \U1/aes_core/SB0/n46 , \U1/aes_core/SB0/n45 ,
         \U1/aes_core/SB0/n44 , \U1/aes_core/SB0/n43 , \U1/aes_core/SB0/n42 ,
         \U1/aes_core/SB0/n41 , \U1/aes_core/SB0/n40 , \U1/aes_core/SB0/n39 ,
         \U1/aes_core/SB0/n38 , \U1/aes_core/SB0/n37 , \U1/aes_core/SB0/n36 ,
         \U1/aes_core/SB0/n35 , \U1/aes_core/SB0/n34 , \U1/aes_core/SB0/n33 ,
         \U1/aes_core/SB0/n32 , \U1/aes_core/SB0/n31 , \U1/aes_core/SB0/n30 ,
         \U1/aes_core/SB0/n29 , \U1/aes_core/SB0/n28 , \U1/aes_core/SB0/n27 ,
         \U1/aes_core/SB0/n26 , \U1/aes_core/SB0/n25 , \U1/aes_core/SB0/n24 ,
         \U1/aes_core/SB0/n23 , \U1/aes_core/SB0/n22 , \U1/aes_core/SB0/n21 ,
         \U1/aes_core/SB0/n20 , \U1/aes_core/SB0/n19 , \U1/aes_core/SB0/n18 ,
         \U1/aes_core/SB0/n17 , \U1/aes_core/SB0/n16 , \U1/aes_core/SB0/n15 ,
         \U1/aes_core/SB0/n14 , \U1/aes_core/SB0/n13 , \U1/aes_core/SB0/n12 ,
         \U1/aes_core/SB0/n11 , \U1/aes_core/SB0/n10 , \U1/aes_core/SB0/n9 ,
         \U1/aes_core/SB0/n8 , \U1/aes_core/SB0/n7 , \U1/aes_core/SB0/n6 ,
         \U1/aes_core/SB0/n5 , \U1/aes_core/SB0/n4 , \U1/aes_core/SB0/n3 ,
         \U1/aes_core/SB0/n2 , \U1/aes_core/SB0/n1 , \U1/aes_core/SB1/n3353 ,
         \U1/aes_core/SB1/n3352 , \U1/aes_core/SB1/n3351 ,
         \U1/aes_core/SB1/n3350 , \U1/aes_core/SB1/n3349 ,
         \U1/aes_core/SB1/n3348 , \U1/aes_core/SB1/n3347 ,
         \U1/aes_core/SB1/n3346 , \U1/aes_core/SB1/n3345 ,
         \U1/aes_core/SB1/n3344 , \U1/aes_core/SB1/n3343 ,
         \U1/aes_core/SB1/n3342 , \U1/aes_core/SB1/n3341 ,
         \U1/aes_core/SB1/n3340 , \U1/aes_core/SB1/n3339 ,
         \U1/aes_core/SB1/n3338 , \U1/aes_core/SB1/n3337 ,
         \U1/aes_core/SB1/n3336 , \U1/aes_core/SB1/n3335 ,
         \U1/aes_core/SB1/n3334 , \U1/aes_core/SB1/n3333 ,
         \U1/aes_core/SB1/n3332 , \U1/aes_core/SB1/n3331 ,
         \U1/aes_core/SB1/n3330 , \U1/aes_core/SB1/n3329 ,
         \U1/aes_core/SB1/n3328 , \U1/aes_core/SB1/n3327 ,
         \U1/aes_core/SB1/n3326 , \U1/aes_core/SB1/n3325 ,
         \U1/aes_core/SB1/n3324 , \U1/aes_core/SB1/n3323 ,
         \U1/aes_core/SB1/n3322 , \U1/aes_core/SB1/n3321 ,
         \U1/aes_core/SB1/n3320 , \U1/aes_core/SB1/n3319 ,
         \U1/aes_core/SB1/n3318 , \U1/aes_core/SB1/n3317 ,
         \U1/aes_core/SB1/n3316 , \U1/aes_core/SB1/n3315 ,
         \U1/aes_core/SB1/n3314 , \U1/aes_core/SB1/n3313 ,
         \U1/aes_core/SB1/n3312 , \U1/aes_core/SB1/n3311 ,
         \U1/aes_core/SB1/n3310 , \U1/aes_core/SB1/n3309 ,
         \U1/aes_core/SB1/n3308 , \U1/aes_core/SB1/n3307 ,
         \U1/aes_core/SB1/n3306 , \U1/aes_core/SB1/n3305 ,
         \U1/aes_core/SB1/n3304 , \U1/aes_core/SB1/n3303 ,
         \U1/aes_core/SB1/n3302 , \U1/aes_core/SB1/n3301 ,
         \U1/aes_core/SB1/n3300 , \U1/aes_core/SB1/n3299 ,
         \U1/aes_core/SB1/n3298 , \U1/aes_core/SB1/n3297 ,
         \U1/aes_core/SB1/n3296 , \U1/aes_core/SB1/n3295 ,
         \U1/aes_core/SB1/n3294 , \U1/aes_core/SB1/n3293 ,
         \U1/aes_core/SB1/n3292 , \U1/aes_core/SB1/n3291 ,
         \U1/aes_core/SB1/n3290 , \U1/aes_core/SB1/n3289 ,
         \U1/aes_core/SB1/n3288 , \U1/aes_core/SB1/n3287 ,
         \U1/aes_core/SB1/n3286 , \U1/aes_core/SB1/n3285 ,
         \U1/aes_core/SB1/n3284 , \U1/aes_core/SB1/n3283 ,
         \U1/aes_core/SB1/n3282 , \U1/aes_core/SB1/n3281 ,
         \U1/aes_core/SB1/n3280 , \U1/aes_core/SB1/n3279 ,
         \U1/aes_core/SB1/n3278 , \U1/aes_core/SB1/n3277 ,
         \U1/aes_core/SB1/n3276 , \U1/aes_core/SB1/n3275 ,
         \U1/aes_core/SB1/n3274 , \U1/aes_core/SB1/n3273 ,
         \U1/aes_core/SB1/n3272 , \U1/aes_core/SB1/n3271 ,
         \U1/aes_core/SB1/n3270 , \U1/aes_core/SB1/n3269 ,
         \U1/aes_core/SB1/n3268 , \U1/aes_core/SB1/n3267 ,
         \U1/aes_core/SB1/n3266 , \U1/aes_core/SB1/n3265 ,
         \U1/aes_core/SB1/n3264 , \U1/aes_core/SB1/n3263 ,
         \U1/aes_core/SB1/n3262 , \U1/aes_core/SB1/n3261 ,
         \U1/aes_core/SB1/n3260 , \U1/aes_core/SB1/n3259 ,
         \U1/aes_core/SB1/n3258 , \U1/aes_core/SB1/n3257 ,
         \U1/aes_core/SB1/n3256 , \U1/aes_core/SB1/n3255 ,
         \U1/aes_core/SB1/n3254 , \U1/aes_core/SB1/n3253 ,
         \U1/aes_core/SB1/n3252 , \U1/aes_core/SB1/n3251 ,
         \U1/aes_core/SB1/n3250 , \U1/aes_core/SB1/n3249 ,
         \U1/aes_core/SB1/n3248 , \U1/aes_core/SB1/n3247 ,
         \U1/aes_core/SB1/n3246 , \U1/aes_core/SB1/n3245 ,
         \U1/aes_core/SB1/n3244 , \U1/aes_core/SB1/n3243 ,
         \U1/aes_core/SB1/n3242 , \U1/aes_core/SB1/n3241 ,
         \U1/aes_core/SB1/n3240 , \U1/aes_core/SB1/n3239 ,
         \U1/aes_core/SB1/n3238 , \U1/aes_core/SB1/n3237 ,
         \U1/aes_core/SB1/n3236 , \U1/aes_core/SB1/n3235 ,
         \U1/aes_core/SB1/n3234 , \U1/aes_core/SB1/n3233 ,
         \U1/aes_core/SB1/n3232 , \U1/aes_core/SB1/n3231 ,
         \U1/aes_core/SB1/n3230 , \U1/aes_core/SB1/n3229 ,
         \U1/aes_core/SB1/n3228 , \U1/aes_core/SB1/n3227 ,
         \U1/aes_core/SB1/n3226 , \U1/aes_core/SB1/n3225 ,
         \U1/aes_core/SB1/n3224 , \U1/aes_core/SB1/n3223 ,
         \U1/aes_core/SB1/n3222 , \U1/aes_core/SB1/n3221 ,
         \U1/aes_core/SB1/n3220 , \U1/aes_core/SB1/n3219 ,
         \U1/aes_core/SB1/n3218 , \U1/aes_core/SB1/n3217 ,
         \U1/aes_core/SB1/n3216 , \U1/aes_core/SB1/n3215 ,
         \U1/aes_core/SB1/n3214 , \U1/aes_core/SB1/n3213 ,
         \U1/aes_core/SB1/n3212 , \U1/aes_core/SB1/n3211 ,
         \U1/aes_core/SB1/n3210 , \U1/aes_core/SB1/n3209 ,
         \U1/aes_core/SB1/n3208 , \U1/aes_core/SB1/n3207 ,
         \U1/aes_core/SB1/n3206 , \U1/aes_core/SB1/n3205 ,
         \U1/aes_core/SB1/n3204 , \U1/aes_core/SB1/n3203 ,
         \U1/aes_core/SB1/n3202 , \U1/aes_core/SB1/n3201 ,
         \U1/aes_core/SB1/n3200 , \U1/aes_core/SB1/n3199 ,
         \U1/aes_core/SB1/n3198 , \U1/aes_core/SB1/n3197 ,
         \U1/aes_core/SB1/n3196 , \U1/aes_core/SB1/n3195 ,
         \U1/aes_core/SB1/n3194 , \U1/aes_core/SB1/n3193 ,
         \U1/aes_core/SB1/n3192 , \U1/aes_core/SB1/n3191 ,
         \U1/aes_core/SB1/n3190 , \U1/aes_core/SB1/n3189 ,
         \U1/aes_core/SB1/n3188 , \U1/aes_core/SB1/n3187 ,
         \U1/aes_core/SB1/n3186 , \U1/aes_core/SB1/n3185 ,
         \U1/aes_core/SB1/n3184 , \U1/aes_core/SB1/n3183 ,
         \U1/aes_core/SB1/n3182 , \U1/aes_core/SB1/n3181 ,
         \U1/aes_core/SB1/n3180 , \U1/aes_core/SB1/n3179 ,
         \U1/aes_core/SB1/n3178 , \U1/aes_core/SB1/n3177 ,
         \U1/aes_core/SB1/n3176 , \U1/aes_core/SB1/n3175 ,
         \U1/aes_core/SB1/n3174 , \U1/aes_core/SB1/n3173 ,
         \U1/aes_core/SB1/n3172 , \U1/aes_core/SB1/n3171 ,
         \U1/aes_core/SB1/n3170 , \U1/aes_core/SB1/n3169 ,
         \U1/aes_core/SB1/n3168 , \U1/aes_core/SB1/n3167 ,
         \U1/aes_core/SB1/n3166 , \U1/aes_core/SB1/n3165 ,
         \U1/aes_core/SB1/n3164 , \U1/aes_core/SB1/n3163 ,
         \U1/aes_core/SB1/n3162 , \U1/aes_core/SB1/n3161 ,
         \U1/aes_core/SB1/n3160 , \U1/aes_core/SB1/n3159 ,
         \U1/aes_core/SB1/n3158 , \U1/aes_core/SB1/n3157 ,
         \U1/aes_core/SB1/n3156 , \U1/aes_core/SB1/n3155 ,
         \U1/aes_core/SB1/n3154 , \U1/aes_core/SB1/n3153 ,
         \U1/aes_core/SB1/n3152 , \U1/aes_core/SB1/n3151 ,
         \U1/aes_core/SB1/n3150 , \U1/aes_core/SB1/n3149 ,
         \U1/aes_core/SB1/n3148 , \U1/aes_core/SB1/n3147 ,
         \U1/aes_core/SB1/n3146 , \U1/aes_core/SB1/n3145 ,
         \U1/aes_core/SB1/n3144 , \U1/aes_core/SB1/n3143 ,
         \U1/aes_core/SB1/n3142 , \U1/aes_core/SB1/n3141 ,
         \U1/aes_core/SB1/n3140 , \U1/aes_core/SB1/n3139 ,
         \U1/aes_core/SB1/n3138 , \U1/aes_core/SB1/n3137 ,
         \U1/aes_core/SB1/n3136 , \U1/aes_core/SB1/n3135 ,
         \U1/aes_core/SB1/n3134 , \U1/aes_core/SB1/n3133 ,
         \U1/aes_core/SB1/n3132 , \U1/aes_core/SB1/n3131 ,
         \U1/aes_core/SB1/n3130 , \U1/aes_core/SB1/n3129 ,
         \U1/aes_core/SB1/n3128 , \U1/aes_core/SB1/n3127 ,
         \U1/aes_core/SB1/n3126 , \U1/aes_core/SB1/n3125 ,
         \U1/aes_core/SB1/n3124 , \U1/aes_core/SB1/n3123 ,
         \U1/aes_core/SB1/n3122 , \U1/aes_core/SB1/n3121 ,
         \U1/aes_core/SB1/n3120 , \U1/aes_core/SB1/n3119 ,
         \U1/aes_core/SB1/n3118 , \U1/aes_core/SB1/n3117 ,
         \U1/aes_core/SB1/n3116 , \U1/aes_core/SB1/n3115 ,
         \U1/aes_core/SB1/n3114 , \U1/aes_core/SB1/n3113 ,
         \U1/aes_core/SB1/n3112 , \U1/aes_core/SB1/n3111 ,
         \U1/aes_core/SB1/n3110 , \U1/aes_core/SB1/n3109 ,
         \U1/aes_core/SB1/n3108 , \U1/aes_core/SB1/n3107 ,
         \U1/aes_core/SB1/n3106 , \U1/aes_core/SB1/n3105 ,
         \U1/aes_core/SB1/n3104 , \U1/aes_core/SB1/n3103 ,
         \U1/aes_core/SB1/n3102 , \U1/aes_core/SB1/n3101 ,
         \U1/aes_core/SB1/n3100 , \U1/aes_core/SB1/n3099 ,
         \U1/aes_core/SB1/n3098 , \U1/aes_core/SB1/n3097 ,
         \U1/aes_core/SB1/n3096 , \U1/aes_core/SB1/n3095 ,
         \U1/aes_core/SB1/n3094 , \U1/aes_core/SB1/n3093 ,
         \U1/aes_core/SB1/n3092 , \U1/aes_core/SB1/n3091 ,
         \U1/aes_core/SB1/n3090 , \U1/aes_core/SB1/n3089 ,
         \U1/aes_core/SB1/n3088 , \U1/aes_core/SB1/n3087 ,
         \U1/aes_core/SB1/n3086 , \U1/aes_core/SB1/n3085 ,
         \U1/aes_core/SB1/n3084 , \U1/aes_core/SB1/n3083 ,
         \U1/aes_core/SB1/n3082 , \U1/aes_core/SB1/n3081 ,
         \U1/aes_core/SB1/n3080 , \U1/aes_core/SB1/n3079 ,
         \U1/aes_core/SB1/n3078 , \U1/aes_core/SB1/n3077 ,
         \U1/aes_core/SB1/n3076 , \U1/aes_core/SB1/n3075 ,
         \U1/aes_core/SB1/n3074 , \U1/aes_core/SB1/n3073 ,
         \U1/aes_core/SB1/n3072 , \U1/aes_core/SB1/n3071 ,
         \U1/aes_core/SB1/n3070 , \U1/aes_core/SB1/n3069 ,
         \U1/aes_core/SB1/n3068 , \U1/aes_core/SB1/n3067 ,
         \U1/aes_core/SB1/n3066 , \U1/aes_core/SB1/n3065 ,
         \U1/aes_core/SB1/n3064 , \U1/aes_core/SB1/n3063 ,
         \U1/aes_core/SB1/n3062 , \U1/aes_core/SB1/n3061 ,
         \U1/aes_core/SB1/n3060 , \U1/aes_core/SB1/n3059 ,
         \U1/aes_core/SB1/n3058 , \U1/aes_core/SB1/n3057 ,
         \U1/aes_core/SB1/n3056 , \U1/aes_core/SB1/n3055 ,
         \U1/aes_core/SB1/n3054 , \U1/aes_core/SB1/n3053 ,
         \U1/aes_core/SB1/n3052 , \U1/aes_core/SB1/n3051 ,
         \U1/aes_core/SB1/n3050 , \U1/aes_core/SB1/n3049 ,
         \U1/aes_core/SB1/n3048 , \U1/aes_core/SB1/n3047 ,
         \U1/aes_core/SB1/n3046 , \U1/aes_core/SB1/n3045 ,
         \U1/aes_core/SB1/n3044 , \U1/aes_core/SB1/n3043 ,
         \U1/aes_core/SB1/n3042 , \U1/aes_core/SB1/n3041 ,
         \U1/aes_core/SB1/n3040 , \U1/aes_core/SB1/n3039 ,
         \U1/aes_core/SB1/n3038 , \U1/aes_core/SB1/n3037 ,
         \U1/aes_core/SB1/n3036 , \U1/aes_core/SB1/n3035 ,
         \U1/aes_core/SB1/n3034 , \U1/aes_core/SB1/n3033 ,
         \U1/aes_core/SB1/n3032 , \U1/aes_core/SB1/n3031 ,
         \U1/aes_core/SB1/n3030 , \U1/aes_core/SB1/n3029 ,
         \U1/aes_core/SB1/n3028 , \U1/aes_core/SB1/n3027 ,
         \U1/aes_core/SB1/n3026 , \U1/aes_core/SB1/n3025 ,
         \U1/aes_core/SB1/n3024 , \U1/aes_core/SB1/n3023 ,
         \U1/aes_core/SB1/n3022 , \U1/aes_core/SB1/n3021 ,
         \U1/aes_core/SB1/n3020 , \U1/aes_core/SB1/n3019 ,
         \U1/aes_core/SB1/n3018 , \U1/aes_core/SB1/n3017 ,
         \U1/aes_core/SB1/n3016 , \U1/aes_core/SB1/n3015 ,
         \U1/aes_core/SB1/n3014 , \U1/aes_core/SB1/n3013 ,
         \U1/aes_core/SB1/n3012 , \U1/aes_core/SB1/n3011 ,
         \U1/aes_core/SB1/n3010 , \U1/aes_core/SB1/n3009 ,
         \U1/aes_core/SB1/n3008 , \U1/aes_core/SB1/n3007 ,
         \U1/aes_core/SB1/n3006 , \U1/aes_core/SB1/n3005 ,
         \U1/aes_core/SB1/n3004 , \U1/aes_core/SB1/n3003 ,
         \U1/aes_core/SB1/n3002 , \U1/aes_core/SB1/n3001 ,
         \U1/aes_core/SB1/n3000 , \U1/aes_core/SB1/n2999 ,
         \U1/aes_core/SB1/n2998 , \U1/aes_core/SB1/n2997 ,
         \U1/aes_core/SB1/n2996 , \U1/aes_core/SB1/n2995 ,
         \U1/aes_core/SB1/n2994 , \U1/aes_core/SB1/n2993 ,
         \U1/aes_core/SB1/n2992 , \U1/aes_core/SB1/n2991 ,
         \U1/aes_core/SB1/n2990 , \U1/aes_core/SB1/n2989 ,
         \U1/aes_core/SB1/n2988 , \U1/aes_core/SB1/n2987 ,
         \U1/aes_core/SB1/n2986 , \U1/aes_core/SB1/n2985 ,
         \U1/aes_core/SB1/n2984 , \U1/aes_core/SB1/n2983 ,
         \U1/aes_core/SB1/n2982 , \U1/aes_core/SB1/n2981 ,
         \U1/aes_core/SB1/n2980 , \U1/aes_core/SB1/n2979 ,
         \U1/aes_core/SB1/n2978 , \U1/aes_core/SB1/n2977 ,
         \U1/aes_core/SB1/n2976 , \U1/aes_core/SB1/n2975 ,
         \U1/aes_core/SB1/n2974 , \U1/aes_core/SB1/n2973 ,
         \U1/aes_core/SB1/n2972 , \U1/aes_core/SB1/n2971 ,
         \U1/aes_core/SB1/n2970 , \U1/aes_core/SB1/n2969 ,
         \U1/aes_core/SB1/n2968 , \U1/aes_core/SB1/n2967 ,
         \U1/aes_core/SB1/n2966 , \U1/aes_core/SB1/n2965 ,
         \U1/aes_core/SB1/n2964 , \U1/aes_core/SB1/n2963 ,
         \U1/aes_core/SB1/n2962 , \U1/aes_core/SB1/n2961 ,
         \U1/aes_core/SB1/n2960 , \U1/aes_core/SB1/n2959 ,
         \U1/aes_core/SB1/n2958 , \U1/aes_core/SB1/n2957 ,
         \U1/aes_core/SB1/n2956 , \U1/aes_core/SB1/n2955 ,
         \U1/aes_core/SB1/n2954 , \U1/aes_core/SB1/n2953 ,
         \U1/aes_core/SB1/n2952 , \U1/aes_core/SB1/n2951 ,
         \U1/aes_core/SB1/n2950 , \U1/aes_core/SB1/n2949 ,
         \U1/aes_core/SB1/n2948 , \U1/aes_core/SB1/n2947 ,
         \U1/aes_core/SB1/n2946 , \U1/aes_core/SB1/n2945 ,
         \U1/aes_core/SB1/n2944 , \U1/aes_core/SB1/n2943 ,
         \U1/aes_core/SB1/n2942 , \U1/aes_core/SB1/n2941 ,
         \U1/aes_core/SB1/n2940 , \U1/aes_core/SB1/n2939 ,
         \U1/aes_core/SB1/n2938 , \U1/aes_core/SB1/n2937 ,
         \U1/aes_core/SB1/n2936 , \U1/aes_core/SB1/n2935 ,
         \U1/aes_core/SB1/n2934 , \U1/aes_core/SB1/n2933 ,
         \U1/aes_core/SB1/n2932 , \U1/aes_core/SB1/n2931 ,
         \U1/aes_core/SB1/n2930 , \U1/aes_core/SB1/n2929 ,
         \U1/aes_core/SB1/n2928 , \U1/aes_core/SB1/n2927 ,
         \U1/aes_core/SB1/n2926 , \U1/aes_core/SB1/n2925 ,
         \U1/aes_core/SB1/n2924 , \U1/aes_core/SB1/n2923 ,
         \U1/aes_core/SB1/n2922 , \U1/aes_core/SB1/n2921 ,
         \U1/aes_core/SB1/n2920 , \U1/aes_core/SB1/n2919 ,
         \U1/aes_core/SB1/n2918 , \U1/aes_core/SB1/n2917 ,
         \U1/aes_core/SB1/n2916 , \U1/aes_core/SB1/n2915 ,
         \U1/aes_core/SB1/n2914 , \U1/aes_core/SB1/n2913 ,
         \U1/aes_core/SB1/n2912 , \U1/aes_core/SB1/n2911 ,
         \U1/aes_core/SB1/n2910 , \U1/aes_core/SB1/n2909 ,
         \U1/aes_core/SB1/n2908 , \U1/aes_core/SB1/n2907 ,
         \U1/aes_core/SB1/n2906 , \U1/aes_core/SB1/n2905 ,
         \U1/aes_core/SB1/n2904 , \U1/aes_core/SB1/n2903 ,
         \U1/aes_core/SB1/n2902 , \U1/aes_core/SB1/n2901 ,
         \U1/aes_core/SB1/n2900 , \U1/aes_core/SB1/n2899 ,
         \U1/aes_core/SB1/n2898 , \U1/aes_core/SB1/n2897 ,
         \U1/aes_core/SB1/n2896 , \U1/aes_core/SB1/n2895 ,
         \U1/aes_core/SB1/n2894 , \U1/aes_core/SB1/n2893 ,
         \U1/aes_core/SB1/n2892 , \U1/aes_core/SB1/n2891 ,
         \U1/aes_core/SB1/n2890 , \U1/aes_core/SB1/n2889 ,
         \U1/aes_core/SB1/n2888 , \U1/aes_core/SB1/n2887 ,
         \U1/aes_core/SB1/n2886 , \U1/aes_core/SB1/n2885 ,
         \U1/aes_core/SB1/n2884 , \U1/aes_core/SB1/n2883 ,
         \U1/aes_core/SB1/n2882 , \U1/aes_core/SB1/n2881 ,
         \U1/aes_core/SB1/n2880 , \U1/aes_core/SB1/n2879 ,
         \U1/aes_core/SB1/n2878 , \U1/aes_core/SB1/n2877 ,
         \U1/aes_core/SB1/n2876 , \U1/aes_core/SB1/n2875 ,
         \U1/aes_core/SB1/n2874 , \U1/aes_core/SB1/n2873 ,
         \U1/aes_core/SB1/n2872 , \U1/aes_core/SB1/n2871 ,
         \U1/aes_core/SB1/n2870 , \U1/aes_core/SB1/n2869 ,
         \U1/aes_core/SB1/n2868 , \U1/aes_core/SB1/n2867 ,
         \U1/aes_core/SB1/n2866 , \U1/aes_core/SB1/n2865 ,
         \U1/aes_core/SB1/n2864 , \U1/aes_core/SB1/n2863 ,
         \U1/aes_core/SB1/n2862 , \U1/aes_core/SB1/n2861 ,
         \U1/aes_core/SB1/n2860 , \U1/aes_core/SB1/n2859 ,
         \U1/aes_core/SB1/n2858 , \U1/aes_core/SB1/n2857 ,
         \U1/aes_core/SB1/n2856 , \U1/aes_core/SB1/n2855 ,
         \U1/aes_core/SB1/n2854 , \U1/aes_core/SB1/n2853 ,
         \U1/aes_core/SB1/n2852 , \U1/aes_core/SB1/n2851 ,
         \U1/aes_core/SB1/n2850 , \U1/aes_core/SB1/n2849 ,
         \U1/aes_core/SB1/n2848 , \U1/aes_core/SB1/n2847 ,
         \U1/aes_core/SB1/n2846 , \U1/aes_core/SB1/n2845 ,
         \U1/aes_core/SB1/n2844 , \U1/aes_core/SB1/n2843 ,
         \U1/aes_core/SB1/n2842 , \U1/aes_core/SB1/n2841 ,
         \U1/aes_core/SB1/n2840 , \U1/aes_core/SB1/n2839 ,
         \U1/aes_core/SB1/n2838 , \U1/aes_core/SB1/n2837 ,
         \U1/aes_core/SB1/n2836 , \U1/aes_core/SB1/n2835 ,
         \U1/aes_core/SB1/n2834 , \U1/aes_core/SB1/n2833 ,
         \U1/aes_core/SB1/n2832 , \U1/aes_core/SB1/n2831 ,
         \U1/aes_core/SB1/n2830 , \U1/aes_core/SB1/n2829 ,
         \U1/aes_core/SB1/n2828 , \U1/aes_core/SB1/n2827 ,
         \U1/aes_core/SB1/n2826 , \U1/aes_core/SB1/n2825 ,
         \U1/aes_core/SB1/n2824 , \U1/aes_core/SB1/n2823 ,
         \U1/aes_core/SB1/n2822 , \U1/aes_core/SB1/n2821 ,
         \U1/aes_core/SB1/n2820 , \U1/aes_core/SB1/n2819 ,
         \U1/aes_core/SB1/n2818 , \U1/aes_core/SB1/n2817 ,
         \U1/aes_core/SB1/n2816 , \U1/aes_core/SB1/n2815 ,
         \U1/aes_core/SB1/n2814 , \U1/aes_core/SB1/n2813 ,
         \U1/aes_core/SB1/n2812 , \U1/aes_core/SB1/n2811 ,
         \U1/aes_core/SB1/n2810 , \U1/aes_core/SB1/n2809 ,
         \U1/aes_core/SB1/n2808 , \U1/aes_core/SB1/n2807 ,
         \U1/aes_core/SB1/n2806 , \U1/aes_core/SB1/n2805 ,
         \U1/aes_core/SB1/n2804 , \U1/aes_core/SB1/n2803 ,
         \U1/aes_core/SB1/n2802 , \U1/aes_core/SB1/n2801 ,
         \U1/aes_core/SB1/n2800 , \U1/aes_core/SB1/n2799 ,
         \U1/aes_core/SB1/n2798 , \U1/aes_core/SB1/n2797 ,
         \U1/aes_core/SB1/n2796 , \U1/aes_core/SB1/n2795 ,
         \U1/aes_core/SB1/n2794 , \U1/aes_core/SB1/n2793 ,
         \U1/aes_core/SB1/n2792 , \U1/aes_core/SB1/n2791 ,
         \U1/aes_core/SB1/n2790 , \U1/aes_core/SB1/n2789 ,
         \U1/aes_core/SB1/n2788 , \U1/aes_core/SB1/n2787 ,
         \U1/aes_core/SB1/n2786 , \U1/aes_core/SB1/n2785 ,
         \U1/aes_core/SB1/n2784 , \U1/aes_core/SB1/n2783 ,
         \U1/aes_core/SB1/n2782 , \U1/aes_core/SB1/n2781 ,
         \U1/aes_core/SB1/n2780 , \U1/aes_core/SB1/n2779 ,
         \U1/aes_core/SB1/n2778 , \U1/aes_core/SB1/n2777 ,
         \U1/aes_core/SB1/n2776 , \U1/aes_core/SB1/n2775 ,
         \U1/aes_core/SB1/n2774 , \U1/aes_core/SB1/n2773 ,
         \U1/aes_core/SB1/n2772 , \U1/aes_core/SB1/n2771 ,
         \U1/aes_core/SB1/n2770 , \U1/aes_core/SB1/n2769 ,
         \U1/aes_core/SB1/n2768 , \U1/aes_core/SB1/n2767 ,
         \U1/aes_core/SB1/n2766 , \U1/aes_core/SB1/n2765 ,
         \U1/aes_core/SB1/n2764 , \U1/aes_core/SB1/n2763 ,
         \U1/aes_core/SB1/n2762 , \U1/aes_core/SB1/n2761 ,
         \U1/aes_core/SB1/n2760 , \U1/aes_core/SB1/n2759 ,
         \U1/aes_core/SB1/n2758 , \U1/aes_core/SB1/n2757 ,
         \U1/aes_core/SB1/n2756 , \U1/aes_core/SB1/n2755 ,
         \U1/aes_core/SB1/n2754 , \U1/aes_core/SB1/n2753 ,
         \U1/aes_core/SB1/n2752 , \U1/aes_core/SB1/n2751 ,
         \U1/aes_core/SB1/n2750 , \U1/aes_core/SB1/n2749 ,
         \U1/aes_core/SB1/n2748 , \U1/aes_core/SB1/n2747 ,
         \U1/aes_core/SB1/n2746 , \U1/aes_core/SB1/n2745 ,
         \U1/aes_core/SB1/n2744 , \U1/aes_core/SB1/n2743 ,
         \U1/aes_core/SB1/n2742 , \U1/aes_core/SB1/n2741 ,
         \U1/aes_core/SB1/n2740 , \U1/aes_core/SB1/n2739 ,
         \U1/aes_core/SB1/n2738 , \U1/aes_core/SB1/n2737 ,
         \U1/aes_core/SB1/n2736 , \U1/aes_core/SB1/n2735 ,
         \U1/aes_core/SB1/n2734 , \U1/aes_core/SB1/n2733 ,
         \U1/aes_core/SB1/n2732 , \U1/aes_core/SB1/n2731 ,
         \U1/aes_core/SB1/n2730 , \U1/aes_core/SB1/n2729 ,
         \U1/aes_core/SB1/n2728 , \U1/aes_core/SB1/n2727 ,
         \U1/aes_core/SB1/n2726 , \U1/aes_core/SB1/n2725 ,
         \U1/aes_core/SB1/n2724 , \U1/aes_core/SB1/n2723 ,
         \U1/aes_core/SB1/n2722 , \U1/aes_core/SB1/n2721 ,
         \U1/aes_core/SB1/n2720 , \U1/aes_core/SB1/n2719 ,
         \U1/aes_core/SB1/n2718 , \U1/aes_core/SB1/n2717 ,
         \U1/aes_core/SB1/n2716 , \U1/aes_core/SB1/n2715 ,
         \U1/aes_core/SB1/n2714 , \U1/aes_core/SB1/n2713 ,
         \U1/aes_core/SB1/n2712 , \U1/aes_core/SB1/n2711 ,
         \U1/aes_core/SB1/n2710 , \U1/aes_core/SB1/n2709 ,
         \U1/aes_core/SB1/n2708 , \U1/aes_core/SB1/n2707 ,
         \U1/aes_core/SB1/n2706 , \U1/aes_core/SB1/n2705 ,
         \U1/aes_core/SB1/n2704 , \U1/aes_core/SB1/n2703 ,
         \U1/aes_core/SB1/n2702 , \U1/aes_core/SB1/n2701 ,
         \U1/aes_core/SB1/n2700 , \U1/aes_core/SB1/n2699 ,
         \U1/aes_core/SB1/n2698 , \U1/aes_core/SB1/n2697 ,
         \U1/aes_core/SB1/n2696 , \U1/aes_core/SB1/n2695 ,
         \U1/aes_core/SB1/n2694 , \U1/aes_core/SB1/n2693 ,
         \U1/aes_core/SB1/n2692 , \U1/aes_core/SB1/n2691 ,
         \U1/aes_core/SB1/n2690 , \U1/aes_core/SB1/n2689 ,
         \U1/aes_core/SB1/n2688 , \U1/aes_core/SB1/n2687 ,
         \U1/aes_core/SB1/n2686 , \U1/aes_core/SB1/n2685 ,
         \U1/aes_core/SB1/n2684 , \U1/aes_core/SB1/n2683 ,
         \U1/aes_core/SB1/n2682 , \U1/aes_core/SB1/n2681 ,
         \U1/aes_core/SB1/n2680 , \U1/aes_core/SB1/n2679 ,
         \U1/aes_core/SB1/n2678 , \U1/aes_core/SB1/n2677 ,
         \U1/aes_core/SB1/n2676 , \U1/aes_core/SB1/n2675 ,
         \U1/aes_core/SB1/n2674 , \U1/aes_core/SB1/n2673 ,
         \U1/aes_core/SB1/n2672 , \U1/aes_core/SB1/n2671 ,
         \U1/aes_core/SB1/n2670 , \U1/aes_core/SB1/n2669 ,
         \U1/aes_core/SB1/n2668 , \U1/aes_core/SB1/n2667 ,
         \U1/aes_core/SB1/n2666 , \U1/aes_core/SB1/n2665 ,
         \U1/aes_core/SB1/n2664 , \U1/aes_core/SB1/n2663 ,
         \U1/aes_core/SB1/n2662 , \U1/aes_core/SB1/n2661 ,
         \U1/aes_core/SB1/n2660 , \U1/aes_core/SB1/n2659 ,
         \U1/aes_core/SB1/n2658 , \U1/aes_core/SB1/n2657 ,
         \U1/aes_core/SB1/n2656 , \U1/aes_core/SB1/n2655 ,
         \U1/aes_core/SB1/n2654 , \U1/aes_core/SB1/n2653 ,
         \U1/aes_core/SB1/n2652 , \U1/aes_core/SB1/n2651 ,
         \U1/aes_core/SB1/n2650 , \U1/aes_core/SB1/n2649 ,
         \U1/aes_core/SB1/n2648 , \U1/aes_core/SB1/n2647 ,
         \U1/aes_core/SB1/n2646 , \U1/aes_core/SB1/n2645 ,
         \U1/aes_core/SB1/n2644 , \U1/aes_core/SB1/n2643 ,
         \U1/aes_core/SB1/n2642 , \U1/aes_core/SB1/n2641 ,
         \U1/aes_core/SB1/n2640 , \U1/aes_core/SB1/n2639 ,
         \U1/aes_core/SB1/n2638 , \U1/aes_core/SB1/n2637 ,
         \U1/aes_core/SB1/n2636 , \U1/aes_core/SB1/n2635 ,
         \U1/aes_core/SB1/n2634 , \U1/aes_core/SB1/n2633 ,
         \U1/aes_core/SB1/n2632 , \U1/aes_core/SB1/n2631 ,
         \U1/aes_core/SB1/n2630 , \U1/aes_core/SB1/n2629 ,
         \U1/aes_core/SB1/n2628 , \U1/aes_core/SB1/n2627 ,
         \U1/aes_core/SB1/n2626 , \U1/aes_core/SB1/n2625 ,
         \U1/aes_core/SB1/n2624 , \U1/aes_core/SB1/n2623 ,
         \U1/aes_core/SB1/n2622 , \U1/aes_core/SB1/n2621 ,
         \U1/aes_core/SB1/n2620 , \U1/aes_core/SB1/n2619 ,
         \U1/aes_core/SB1/n2618 , \U1/aes_core/SB1/n2617 ,
         \U1/aes_core/SB1/n2616 , \U1/aes_core/SB1/n2615 ,
         \U1/aes_core/SB1/n2614 , \U1/aes_core/SB1/n2613 ,
         \U1/aes_core/SB1/n2612 , \U1/aes_core/SB1/n2611 ,
         \U1/aes_core/SB1/n2610 , \U1/aes_core/SB1/n2609 ,
         \U1/aes_core/SB1/n2608 , \U1/aes_core/SB1/n2607 ,
         \U1/aes_core/SB1/n2606 , \U1/aes_core/SB1/n2605 ,
         \U1/aes_core/SB1/n2604 , \U1/aes_core/SB1/n2603 ,
         \U1/aes_core/SB1/n2602 , \U1/aes_core/SB1/n2601 ,
         \U1/aes_core/SB1/n2600 , \U1/aes_core/SB1/n2599 ,
         \U1/aes_core/SB1/n2598 , \U1/aes_core/SB1/n2597 ,
         \U1/aes_core/SB1/n2596 , \U1/aes_core/SB1/n2595 ,
         \U1/aes_core/SB1/n2594 , \U1/aes_core/SB1/n2593 ,
         \U1/aes_core/SB1/n2592 , \U1/aes_core/SB1/n2591 ,
         \U1/aes_core/SB1/n2590 , \U1/aes_core/SB1/n2589 ,
         \U1/aes_core/SB1/n2588 , \U1/aes_core/SB1/n2587 ,
         \U1/aes_core/SB1/n2586 , \U1/aes_core/SB1/n2585 ,
         \U1/aes_core/SB1/n2584 , \U1/aes_core/SB1/n2583 ,
         \U1/aes_core/SB1/n2582 , \U1/aes_core/SB1/n2581 ,
         \U1/aes_core/SB1/n2580 , \U1/aes_core/SB1/n2579 ,
         \U1/aes_core/SB1/n2578 , \U1/aes_core/SB1/n2577 ,
         \U1/aes_core/SB1/n2576 , \U1/aes_core/SB1/n2575 ,
         \U1/aes_core/SB1/n2574 , \U1/aes_core/SB1/n2573 ,
         \U1/aes_core/SB1/n2572 , \U1/aes_core/SB1/n2571 ,
         \U1/aes_core/SB1/n2570 , \U1/aes_core/SB1/n2569 ,
         \U1/aes_core/SB1/n2568 , \U1/aes_core/SB1/n2567 ,
         \U1/aes_core/SB1/n2566 , \U1/aes_core/SB1/n2565 ,
         \U1/aes_core/SB1/n2564 , \U1/aes_core/SB1/n2563 ,
         \U1/aes_core/SB1/n2562 , \U1/aes_core/SB1/n2561 ,
         \U1/aes_core/SB1/n2560 , \U1/aes_core/SB1/n2559 ,
         \U1/aes_core/SB1/n2558 , \U1/aes_core/SB1/n2557 ,
         \U1/aes_core/SB1/n2556 , \U1/aes_core/SB1/n2555 ,
         \U1/aes_core/SB1/n2554 , \U1/aes_core/SB1/n2553 ,
         \U1/aes_core/SB1/n2552 , \U1/aes_core/SB1/n2551 ,
         \U1/aes_core/SB1/n2550 , \U1/aes_core/SB1/n2549 ,
         \U1/aes_core/SB1/n2548 , \U1/aes_core/SB1/n2547 ,
         \U1/aes_core/SB1/n2546 , \U1/aes_core/SB1/n2545 ,
         \U1/aes_core/SB1/n2544 , \U1/aes_core/SB1/n2543 ,
         \U1/aes_core/SB1/n2542 , \U1/aes_core/SB1/n2541 ,
         \U1/aes_core/SB1/n2540 , \U1/aes_core/SB1/n2539 ,
         \U1/aes_core/SB1/n2538 , \U1/aes_core/SB1/n2537 ,
         \U1/aes_core/SB1/n2536 , \U1/aes_core/SB1/n2535 ,
         \U1/aes_core/SB1/n2534 , \U1/aes_core/SB1/n2533 ,
         \U1/aes_core/SB1/n2532 , \U1/aes_core/SB1/n2531 ,
         \U1/aes_core/SB1/n2530 , \U1/aes_core/SB1/n2529 ,
         \U1/aes_core/SB1/n2528 , \U1/aes_core/SB1/n2527 ,
         \U1/aes_core/SB1/n2526 , \U1/aes_core/SB1/n2525 ,
         \U1/aes_core/SB1/n2524 , \U1/aes_core/SB1/n2523 ,
         \U1/aes_core/SB1/n2522 , \U1/aes_core/SB1/n2521 ,
         \U1/aes_core/SB1/n2520 , \U1/aes_core/SB1/n2519 ,
         \U1/aes_core/SB1/n2518 , \U1/aes_core/SB1/n2517 ,
         \U1/aes_core/SB1/n2516 , \U1/aes_core/SB1/n2515 ,
         \U1/aes_core/SB1/n2514 , \U1/aes_core/SB1/n2513 ,
         \U1/aes_core/SB1/n2512 , \U1/aes_core/SB1/n2511 ,
         \U1/aes_core/SB1/n2510 , \U1/aes_core/SB1/n2509 ,
         \U1/aes_core/SB1/n2508 , \U1/aes_core/SB1/n2507 ,
         \U1/aes_core/SB1/n2506 , \U1/aes_core/SB1/n2505 ,
         \U1/aes_core/SB1/n2504 , \U1/aes_core/SB1/n2503 ,
         \U1/aes_core/SB1/n2502 , \U1/aes_core/SB1/n2501 ,
         \U1/aes_core/SB1/n2500 , \U1/aes_core/SB1/n2499 ,
         \U1/aes_core/SB1/n2498 , \U1/aes_core/SB1/n2497 ,
         \U1/aes_core/SB1/n2496 , \U1/aes_core/SB1/n2495 ,
         \U1/aes_core/SB1/n2494 , \U1/aes_core/SB1/n2493 ,
         \U1/aes_core/SB1/n2492 , \U1/aes_core/SB1/n2491 ,
         \U1/aes_core/SB1/n2490 , \U1/aes_core/SB1/n2489 ,
         \U1/aes_core/SB1/n2488 , \U1/aes_core/SB1/n2487 ,
         \U1/aes_core/SB1/n2486 , \U1/aes_core/SB1/n2485 ,
         \U1/aes_core/SB1/n2484 , \U1/aes_core/SB1/n2483 ,
         \U1/aes_core/SB1/n2482 , \U1/aes_core/SB1/n2481 ,
         \U1/aes_core/SB1/n2480 , \U1/aes_core/SB1/n2479 ,
         \U1/aes_core/SB1/n2478 , \U1/aes_core/SB1/n2477 ,
         \U1/aes_core/SB1/n2476 , \U1/aes_core/SB1/n2475 ,
         \U1/aes_core/SB1/n2474 , \U1/aes_core/SB1/n2473 ,
         \U1/aes_core/SB1/n2472 , \U1/aes_core/SB1/n2471 ,
         \U1/aes_core/SB1/n2470 , \U1/aes_core/SB1/n2469 ,
         \U1/aes_core/SB1/n2468 , \U1/aes_core/SB1/n2467 ,
         \U1/aes_core/SB1/n2466 , \U1/aes_core/SB1/n2465 ,
         \U1/aes_core/SB1/n2464 , \U1/aes_core/SB1/n2463 ,
         \U1/aes_core/SB1/n2462 , \U1/aes_core/SB1/n2461 ,
         \U1/aes_core/SB1/n2460 , \U1/aes_core/SB1/n2459 ,
         \U1/aes_core/SB1/n2458 , \U1/aes_core/SB1/n2457 ,
         \U1/aes_core/SB1/n2456 , \U1/aes_core/SB1/n2455 ,
         \U1/aes_core/SB1/n2454 , \U1/aes_core/SB1/n2453 ,
         \U1/aes_core/SB1/n2452 , \U1/aes_core/SB1/n2451 ,
         \U1/aes_core/SB1/n2450 , \U1/aes_core/SB1/n2449 ,
         \U1/aes_core/SB1/n2448 , \U1/aes_core/SB1/n2447 ,
         \U1/aes_core/SB1/n2446 , \U1/aes_core/SB1/n2445 ,
         \U1/aes_core/SB1/n2444 , \U1/aes_core/SB1/n2443 ,
         \U1/aes_core/SB1/n2442 , \U1/aes_core/SB1/n2441 ,
         \U1/aes_core/SB1/n2440 , \U1/aes_core/SB1/n2439 ,
         \U1/aes_core/SB1/n2438 , \U1/aes_core/SB1/n2437 ,
         \U1/aes_core/SB1/n2436 , \U1/aes_core/SB1/n2435 ,
         \U1/aes_core/SB1/n2434 , \U1/aes_core/SB1/n2433 ,
         \U1/aes_core/SB1/n2432 , \U1/aes_core/SB1/n2431 ,
         \U1/aes_core/SB1/n2430 , \U1/aes_core/SB1/n2429 ,
         \U1/aes_core/SB1/n2428 , \U1/aes_core/SB1/n2427 ,
         \U1/aes_core/SB1/n2426 , \U1/aes_core/SB1/n2425 ,
         \U1/aes_core/SB1/n2424 , \U1/aes_core/SB1/n2423 ,
         \U1/aes_core/SB1/n2422 , \U1/aes_core/SB1/n2421 ,
         \U1/aes_core/SB1/n2420 , \U1/aes_core/SB1/n2419 ,
         \U1/aes_core/SB1/n2418 , \U1/aes_core/SB1/n2417 ,
         \U1/aes_core/SB1/n2416 , \U1/aes_core/SB1/n2415 ,
         \U1/aes_core/SB1/n2414 , \U1/aes_core/SB1/n2413 ,
         \U1/aes_core/SB1/n2412 , \U1/aes_core/SB1/n2411 ,
         \U1/aes_core/SB1/n2410 , \U1/aes_core/SB1/n2409 ,
         \U1/aes_core/SB1/n2408 , \U1/aes_core/SB1/n2407 ,
         \U1/aes_core/SB1/n2406 , \U1/aes_core/SB1/n2405 ,
         \U1/aes_core/SB1/n2404 , \U1/aes_core/SB1/n2403 ,
         \U1/aes_core/SB1/n2402 , \U1/aes_core/SB1/n2401 ,
         \U1/aes_core/SB1/n2400 , \U1/aes_core/SB1/n2399 ,
         \U1/aes_core/SB1/n2398 , \U1/aes_core/SB1/n2397 ,
         \U1/aes_core/SB1/n2396 , \U1/aes_core/SB1/n2395 ,
         \U1/aes_core/SB1/n2394 , \U1/aes_core/SB1/n2393 ,
         \U1/aes_core/SB1/n2392 , \U1/aes_core/SB1/n2391 ,
         \U1/aes_core/SB1/n2390 , \U1/aes_core/SB1/n2389 ,
         \U1/aes_core/SB1/n2388 , \U1/aes_core/SB1/n2387 ,
         \U1/aes_core/SB1/n2386 , \U1/aes_core/SB1/n2385 ,
         \U1/aes_core/SB1/n2384 , \U1/aes_core/SB1/n2383 ,
         \U1/aes_core/SB1/n2382 , \U1/aes_core/SB1/n2381 ,
         \U1/aes_core/SB1/n2380 , \U1/aes_core/SB1/n2379 ,
         \U1/aes_core/SB1/n2378 , \U1/aes_core/SB1/n2377 ,
         \U1/aes_core/SB1/n2376 , \U1/aes_core/SB1/n2375 ,
         \U1/aes_core/SB1/n2374 , \U1/aes_core/SB1/n2373 ,
         \U1/aes_core/SB1/n2372 , \U1/aes_core/SB1/n2371 ,
         \U1/aes_core/SB1/n2370 , \U1/aes_core/SB1/n2369 ,
         \U1/aes_core/SB1/n2368 , \U1/aes_core/SB1/n2367 ,
         \U1/aes_core/SB1/n2366 , \U1/aes_core/SB1/n2365 ,
         \U1/aes_core/SB1/n2364 , \U1/aes_core/SB1/n2363 ,
         \U1/aes_core/SB1/n2362 , \U1/aes_core/SB1/n2361 ,
         \U1/aes_core/SB1/n2360 , \U1/aes_core/SB1/n2359 ,
         \U1/aes_core/SB1/n2358 , \U1/aes_core/SB1/n2357 ,
         \U1/aes_core/SB1/n2356 , \U1/aes_core/SB1/n2355 ,
         \U1/aes_core/SB1/n2354 , \U1/aes_core/SB1/n2353 ,
         \U1/aes_core/SB1/n2352 , \U1/aes_core/SB1/n2351 ,
         \U1/aes_core/SB1/n2350 , \U1/aes_core/SB1/n2349 ,
         \U1/aes_core/SB1/n2348 , \U1/aes_core/SB1/n2347 ,
         \U1/aes_core/SB1/n2346 , \U1/aes_core/SB1/n2345 ,
         \U1/aes_core/SB1/n2344 , \U1/aes_core/SB1/n2343 ,
         \U1/aes_core/SB1/n2342 , \U1/aes_core/SB1/n2341 ,
         \U1/aes_core/SB1/n2340 , \U1/aes_core/SB1/n2339 ,
         \U1/aes_core/SB1/n2338 , \U1/aes_core/SB1/n2337 ,
         \U1/aes_core/SB1/n2336 , \U1/aes_core/SB1/n2335 ,
         \U1/aes_core/SB1/n2334 , \U1/aes_core/SB1/n2333 ,
         \U1/aes_core/SB1/n2332 , \U1/aes_core/SB1/n2331 ,
         \U1/aes_core/SB1/n2330 , \U1/aes_core/SB1/n2329 ,
         \U1/aes_core/SB1/n2328 , \U1/aes_core/SB1/n2327 ,
         \U1/aes_core/SB1/n2326 , \U1/aes_core/SB1/n2325 ,
         \U1/aes_core/SB1/n2324 , \U1/aes_core/SB1/n2323 ,
         \U1/aes_core/SB1/n2322 , \U1/aes_core/SB1/n2321 ,
         \U1/aes_core/SB1/n2320 , \U1/aes_core/SB1/n2319 ,
         \U1/aes_core/SB1/n2318 , \U1/aes_core/SB1/n2317 ,
         \U1/aes_core/SB1/n2316 , \U1/aes_core/SB1/n2315 ,
         \U1/aes_core/SB1/n2314 , \U1/aes_core/SB1/n2313 ,
         \U1/aes_core/SB1/n2312 , \U1/aes_core/SB1/n2311 ,
         \U1/aes_core/SB1/n2310 , \U1/aes_core/SB1/n2309 ,
         \U1/aes_core/SB1/n2308 , \U1/aes_core/SB1/n2307 ,
         \U1/aes_core/SB1/n2306 , \U1/aes_core/SB1/n2305 ,
         \U1/aes_core/SB1/n2304 , \U1/aes_core/SB1/n2303 ,
         \U1/aes_core/SB1/n2302 , \U1/aes_core/SB1/n2301 ,
         \U1/aes_core/SB1/n2300 , \U1/aes_core/SB1/n2299 ,
         \U1/aes_core/SB1/n2298 , \U1/aes_core/SB1/n2297 ,
         \U1/aes_core/SB1/n2296 , \U1/aes_core/SB1/n2295 ,
         \U1/aes_core/SB1/n2294 , \U1/aes_core/SB1/n2293 ,
         \U1/aes_core/SB1/n2292 , \U1/aes_core/SB1/n2291 ,
         \U1/aes_core/SB1/n2290 , \U1/aes_core/SB1/n2289 ,
         \U1/aes_core/SB1/n2288 , \U1/aes_core/SB1/n2287 ,
         \U1/aes_core/SB1/n2286 , \U1/aes_core/SB1/n2285 ,
         \U1/aes_core/SB1/n2284 , \U1/aes_core/SB1/n2283 ,
         \U1/aes_core/SB1/n2282 , \U1/aes_core/SB1/n2281 ,
         \U1/aes_core/SB1/n2280 , \U1/aes_core/SB1/n2279 ,
         \U1/aes_core/SB1/n2278 , \U1/aes_core/SB1/n2277 ,
         \U1/aes_core/SB1/n2276 , \U1/aes_core/SB1/n2275 ,
         \U1/aes_core/SB1/n2274 , \U1/aes_core/SB1/n2273 ,
         \U1/aes_core/SB1/n2272 , \U1/aes_core/SB1/n2271 ,
         \U1/aes_core/SB1/n2270 , \U1/aes_core/SB1/n2269 ,
         \U1/aes_core/SB1/n2268 , \U1/aes_core/SB1/n2267 ,
         \U1/aes_core/SB1/n2266 , \U1/aes_core/SB1/n2265 ,
         \U1/aes_core/SB1/n2264 , \U1/aes_core/SB1/n2263 ,
         \U1/aes_core/SB1/n2262 , \U1/aes_core/SB1/n2261 ,
         \U1/aes_core/SB1/n2260 , \U1/aes_core/SB1/n2259 ,
         \U1/aes_core/SB1/n2258 , \U1/aes_core/SB1/n2257 ,
         \U1/aes_core/SB1/n2256 , \U1/aes_core/SB1/n2255 ,
         \U1/aes_core/SB1/n2254 , \U1/aes_core/SB1/n2253 ,
         \U1/aes_core/SB1/n2252 , \U1/aes_core/SB1/n2251 ,
         \U1/aes_core/SB1/n2250 , \U1/aes_core/SB1/n2249 ,
         \U1/aes_core/SB1/n2248 , \U1/aes_core/SB1/n2247 ,
         \U1/aes_core/SB1/n2246 , \U1/aes_core/SB1/n2245 ,
         \U1/aes_core/SB1/n2244 , \U1/aes_core/SB1/n2243 ,
         \U1/aes_core/SB1/n2242 , \U1/aes_core/SB1/n2241 ,
         \U1/aes_core/SB1/n2240 , \U1/aes_core/SB1/n2239 ,
         \U1/aes_core/SB1/n2238 , \U1/aes_core/SB1/n2237 ,
         \U1/aes_core/SB1/n2236 , \U1/aes_core/SB1/n2235 ,
         \U1/aes_core/SB1/n2234 , \U1/aes_core/SB1/n2233 ,
         \U1/aes_core/SB1/n2232 , \U1/aes_core/SB1/n2231 ,
         \U1/aes_core/SB1/n2230 , \U1/aes_core/SB1/n2229 ,
         \U1/aes_core/SB1/n2228 , \U1/aes_core/SB1/n2227 ,
         \U1/aes_core/SB1/n2226 , \U1/aes_core/SB1/n2225 ,
         \U1/aes_core/SB1/n2224 , \U1/aes_core/SB1/n2223 ,
         \U1/aes_core/SB1/n2222 , \U1/aes_core/SB1/n2221 ,
         \U1/aes_core/SB1/n2220 , \U1/aes_core/SB1/n2219 ,
         \U1/aes_core/SB1/n2218 , \U1/aes_core/SB1/n2217 ,
         \U1/aes_core/SB1/n2216 , \U1/aes_core/SB1/n2215 ,
         \U1/aes_core/SB1/n2214 , \U1/aes_core/SB1/n2213 ,
         \U1/aes_core/SB1/n2212 , \U1/aes_core/SB1/n2211 ,
         \U1/aes_core/SB1/n2210 , \U1/aes_core/SB1/n2209 ,
         \U1/aes_core/SB1/n2208 , \U1/aes_core/SB1/n2207 ,
         \U1/aes_core/SB1/n2206 , \U1/aes_core/SB1/n2205 ,
         \U1/aes_core/SB1/n2204 , \U1/aes_core/SB1/n2203 ,
         \U1/aes_core/SB1/n2202 , \U1/aes_core/SB1/n2201 ,
         \U1/aes_core/SB1/n2200 , \U1/aes_core/SB1/n2199 ,
         \U1/aes_core/SB1/n2198 , \U1/aes_core/SB1/n2197 ,
         \U1/aes_core/SB1/n2196 , \U1/aes_core/SB1/n2195 ,
         \U1/aes_core/SB1/n2194 , \U1/aes_core/SB1/n2193 ,
         \U1/aes_core/SB1/n2192 , \U1/aes_core/SB1/n2191 ,
         \U1/aes_core/SB1/n2190 , \U1/aes_core/SB1/n2189 ,
         \U1/aes_core/SB1/n2188 , \U1/aes_core/SB1/n2187 ,
         \U1/aes_core/SB1/n2186 , \U1/aes_core/SB1/n2185 ,
         \U1/aes_core/SB1/n2184 , \U1/aes_core/SB1/n2183 ,
         \U1/aes_core/SB1/n2182 , \U1/aes_core/SB1/n2181 ,
         \U1/aes_core/SB1/n2180 , \U1/aes_core/SB1/n2179 ,
         \U1/aes_core/SB1/n2178 , \U1/aes_core/SB1/n2177 ,
         \U1/aes_core/SB1/n2176 , \U1/aes_core/SB1/n2175 ,
         \U1/aes_core/SB1/n2174 , \U1/aes_core/SB1/n2173 ,
         \U1/aes_core/SB1/n2172 , \U1/aes_core/SB1/n2171 ,
         \U1/aes_core/SB1/n2170 , \U1/aes_core/SB1/n2169 ,
         \U1/aes_core/SB1/n2168 , \U1/aes_core/SB1/n2167 ,
         \U1/aes_core/SB1/n2166 , \U1/aes_core/SB1/n2165 ,
         \U1/aes_core/SB1/n2164 , \U1/aes_core/SB1/n2163 ,
         \U1/aes_core/SB1/n2162 , \U1/aes_core/SB1/n2161 ,
         \U1/aes_core/SB1/n2160 , \U1/aes_core/SB1/n2159 ,
         \U1/aes_core/SB1/n2158 , \U1/aes_core/SB1/n2157 ,
         \U1/aes_core/SB1/n2156 , \U1/aes_core/SB1/n2155 ,
         \U1/aes_core/SB1/n2154 , \U1/aes_core/SB1/n2153 ,
         \U1/aes_core/SB1/n2152 , \U1/aes_core/SB1/n2151 ,
         \U1/aes_core/SB1/n2150 , \U1/aes_core/SB1/n2149 ,
         \U1/aes_core/SB1/n2148 , \U1/aes_core/SB1/n2147 ,
         \U1/aes_core/SB1/n2146 , \U1/aes_core/SB1/n2145 ,
         \U1/aes_core/SB1/n2144 , \U1/aes_core/SB1/n2143 ,
         \U1/aes_core/SB1/n2142 , \U1/aes_core/SB1/n2141 ,
         \U1/aes_core/SB1/n2140 , \U1/aes_core/SB1/n2139 ,
         \U1/aes_core/SB1/n2138 , \U1/aes_core/SB1/n2137 ,
         \U1/aes_core/SB1/n2136 , \U1/aes_core/SB1/n2135 ,
         \U1/aes_core/SB1/n2134 , \U1/aes_core/SB1/n2133 ,
         \U1/aes_core/SB1/n2132 , \U1/aes_core/SB1/n2131 ,
         \U1/aes_core/SB1/n2130 , \U1/aes_core/SB1/n2129 ,
         \U1/aes_core/SB1/n2128 , \U1/aes_core/SB1/n2127 ,
         \U1/aes_core/SB1/n2126 , \U1/aes_core/SB1/n2125 ,
         \U1/aes_core/SB1/n2124 , \U1/aes_core/SB1/n2123 ,
         \U1/aes_core/SB1/n2122 , \U1/aes_core/SB1/n2121 ,
         \U1/aes_core/SB1/n2120 , \U1/aes_core/SB1/n2119 ,
         \U1/aes_core/SB1/n2118 , \U1/aes_core/SB1/n2117 ,
         \U1/aes_core/SB1/n2116 , \U1/aes_core/SB1/n2115 ,
         \U1/aes_core/SB1/n2114 , \U1/aes_core/SB1/n2113 ,
         \U1/aes_core/SB1/n2112 , \U1/aes_core/SB1/n2111 ,
         \U1/aes_core/SB1/n2110 , \U1/aes_core/SB1/n2109 ,
         \U1/aes_core/SB1/n2108 , \U1/aes_core/SB1/n2107 ,
         \U1/aes_core/SB1/n2106 , \U1/aes_core/SB1/n2105 ,
         \U1/aes_core/SB1/n2104 , \U1/aes_core/SB1/n2103 ,
         \U1/aes_core/SB1/n2102 , \U1/aes_core/SB1/n2101 ,
         \U1/aes_core/SB1/n2100 , \U1/aes_core/SB1/n2099 ,
         \U1/aes_core/SB1/n2098 , \U1/aes_core/SB1/n2097 ,
         \U1/aes_core/SB1/n2096 , \U1/aes_core/SB1/n2095 ,
         \U1/aes_core/SB1/n2094 , \U1/aes_core/SB1/n2093 ,
         \U1/aes_core/SB1/n2092 , \U1/aes_core/SB1/n2091 ,
         \U1/aes_core/SB1/n2090 , \U1/aes_core/SB1/n2089 ,
         \U1/aes_core/SB1/n2088 , \U1/aes_core/SB1/n2087 ,
         \U1/aes_core/SB1/n2086 , \U1/aes_core/SB1/n2085 ,
         \U1/aes_core/SB1/n2084 , \U1/aes_core/SB1/n2083 ,
         \U1/aes_core/SB1/n2082 , \U1/aes_core/SB1/n2081 ,
         \U1/aes_core/SB1/n2080 , \U1/aes_core/SB1/n2079 ,
         \U1/aes_core/SB1/n2078 , \U1/aes_core/SB1/n2077 ,
         \U1/aes_core/SB1/n2076 , \U1/aes_core/SB1/n2075 ,
         \U1/aes_core/SB1/n2074 , \U1/aes_core/SB1/n2073 ,
         \U1/aes_core/SB1/n2072 , \U1/aes_core/SB1/n2071 ,
         \U1/aes_core/SB1/n2070 , \U1/aes_core/SB1/n2069 ,
         \U1/aes_core/SB1/n2068 , \U1/aes_core/SB1/n2067 ,
         \U1/aes_core/SB1/n2066 , \U1/aes_core/SB1/n2065 ,
         \U1/aes_core/SB1/n2064 , \U1/aes_core/SB1/n2063 ,
         \U1/aes_core/SB1/n2062 , \U1/aes_core/SB1/n2061 ,
         \U1/aes_core/SB1/n2060 , \U1/aes_core/SB1/n2059 ,
         \U1/aes_core/SB1/n2058 , \U1/aes_core/SB1/n2057 ,
         \U1/aes_core/SB1/n2056 , \U1/aes_core/SB1/n2055 ,
         \U1/aes_core/SB1/n2054 , \U1/aes_core/SB1/n2053 ,
         \U1/aes_core/SB1/n2052 , \U1/aes_core/SB1/n2051 ,
         \U1/aes_core/SB1/n2050 , \U1/aes_core/SB1/n2049 ,
         \U1/aes_core/SB1/n2048 , \U1/aes_core/SB1/n2047 ,
         \U1/aes_core/SB1/n2046 , \U1/aes_core/SB1/n2045 ,
         \U1/aes_core/SB1/n2044 , \U1/aes_core/SB1/n2043 ,
         \U1/aes_core/SB1/n2042 , \U1/aes_core/SB1/n2041 ,
         \U1/aes_core/SB1/n2040 , \U1/aes_core/SB1/n2039 ,
         \U1/aes_core/SB1/n2038 , \U1/aes_core/SB1/n2037 ,
         \U1/aes_core/SB1/n2036 , \U1/aes_core/SB1/n2035 ,
         \U1/aes_core/SB1/n2034 , \U1/aes_core/SB1/n2033 ,
         \U1/aes_core/SB1/n2032 , \U1/aes_core/SB1/n2031 ,
         \U1/aes_core/SB1/n2030 , \U1/aes_core/SB1/n2029 ,
         \U1/aes_core/SB1/n2028 , \U1/aes_core/SB1/n2027 ,
         \U1/aes_core/SB1/n2026 , \U1/aes_core/SB1/n2025 ,
         \U1/aes_core/SB1/n2024 , \U1/aes_core/SB1/n2023 ,
         \U1/aes_core/SB1/n2022 , \U1/aes_core/SB1/n2021 ,
         \U1/aes_core/SB1/n2020 , \U1/aes_core/SB1/n2019 ,
         \U1/aes_core/SB1/n2018 , \U1/aes_core/SB1/n2017 ,
         \U1/aes_core/SB1/n2016 , \U1/aes_core/SB1/n2015 ,
         \U1/aes_core/SB1/n2014 , \U1/aes_core/SB1/n2013 ,
         \U1/aes_core/SB1/n2012 , \U1/aes_core/SB1/n2011 ,
         \U1/aes_core/SB1/n2010 , \U1/aes_core/SB1/n2009 ,
         \U1/aes_core/SB1/n2008 , \U1/aes_core/SB1/n2007 ,
         \U1/aes_core/SB1/n2006 , \U1/aes_core/SB1/n2005 ,
         \U1/aes_core/SB1/n2004 , \U1/aes_core/SB1/n2003 ,
         \U1/aes_core/SB1/n2002 , \U1/aes_core/SB1/n2001 ,
         \U1/aes_core/SB1/n2000 , \U1/aes_core/SB1/n1999 ,
         \U1/aes_core/SB1/n1998 , \U1/aes_core/SB1/n1997 ,
         \U1/aes_core/SB1/n1996 , \U1/aes_core/SB1/n1995 ,
         \U1/aes_core/SB1/n1994 , \U1/aes_core/SB1/n1993 ,
         \U1/aes_core/SB1/n1992 , \U1/aes_core/SB1/n1991 ,
         \U1/aes_core/SB1/n1990 , \U1/aes_core/SB1/n1989 ,
         \U1/aes_core/SB1/n1988 , \U1/aes_core/SB1/n1987 ,
         \U1/aes_core/SB1/n1986 , \U1/aes_core/SB1/n1985 ,
         \U1/aes_core/SB1/n1984 , \U1/aes_core/SB1/n1983 ,
         \U1/aes_core/SB1/n1982 , \U1/aes_core/SB1/n1981 ,
         \U1/aes_core/SB1/n1980 , \U1/aes_core/SB1/n1979 ,
         \U1/aes_core/SB1/n1978 , \U1/aes_core/SB1/n1977 ,
         \U1/aes_core/SB1/n1976 , \U1/aes_core/SB1/n1975 ,
         \U1/aes_core/SB1/n1974 , \U1/aes_core/SB1/n1973 ,
         \U1/aes_core/SB1/n1972 , \U1/aes_core/SB1/n1971 ,
         \U1/aes_core/SB1/n1970 , \U1/aes_core/SB1/n1969 ,
         \U1/aes_core/SB1/n1968 , \U1/aes_core/SB1/n1967 ,
         \U1/aes_core/SB1/n1966 , \U1/aes_core/SB1/n1965 ,
         \U1/aes_core/SB1/n1964 , \U1/aes_core/SB1/n1963 ,
         \U1/aes_core/SB1/n1962 , \U1/aes_core/SB1/n1961 ,
         \U1/aes_core/SB1/n1960 , \U1/aes_core/SB1/n1959 ,
         \U1/aes_core/SB1/n1958 , \U1/aes_core/SB1/n1957 ,
         \U1/aes_core/SB1/n1956 , \U1/aes_core/SB1/n1955 ,
         \U1/aes_core/SB1/n1954 , \U1/aes_core/SB1/n1953 ,
         \U1/aes_core/SB1/n1952 , \U1/aes_core/SB1/n1951 ,
         \U1/aes_core/SB1/n1950 , \U1/aes_core/SB1/n1949 ,
         \U1/aes_core/SB1/n1948 , \U1/aes_core/SB1/n1947 ,
         \U1/aes_core/SB1/n1946 , \U1/aes_core/SB1/n1945 ,
         \U1/aes_core/SB1/n1944 , \U1/aes_core/SB1/n1943 ,
         \U1/aes_core/SB1/n1942 , \U1/aes_core/SB1/n1941 ,
         \U1/aes_core/SB1/n1940 , \U1/aes_core/SB1/n1939 ,
         \U1/aes_core/SB1/n1938 , \U1/aes_core/SB1/n1937 ,
         \U1/aes_core/SB1/n1936 , \U1/aes_core/SB1/n1935 ,
         \U1/aes_core/SB1/n1934 , \U1/aes_core/SB1/n1933 ,
         \U1/aes_core/SB1/n1932 , \U1/aes_core/SB1/n1931 ,
         \U1/aes_core/SB1/n1930 , \U1/aes_core/SB1/n1929 ,
         \U1/aes_core/SB1/n1928 , \U1/aes_core/SB1/n1927 ,
         \U1/aes_core/SB1/n1926 , \U1/aes_core/SB1/n1925 ,
         \U1/aes_core/SB1/n1924 , \U1/aes_core/SB1/n1923 ,
         \U1/aes_core/SB1/n1922 , \U1/aes_core/SB1/n1921 ,
         \U1/aes_core/SB1/n1920 , \U1/aes_core/SB1/n1919 ,
         \U1/aes_core/SB1/n1918 , \U1/aes_core/SB1/n1917 ,
         \U1/aes_core/SB1/n1916 , \U1/aes_core/SB1/n1915 ,
         \U1/aes_core/SB1/n1914 , \U1/aes_core/SB1/n1913 ,
         \U1/aes_core/SB1/n1912 , \U1/aes_core/SB1/n1911 ,
         \U1/aes_core/SB1/n1910 , \U1/aes_core/SB1/n1909 ,
         \U1/aes_core/SB1/n1908 , \U1/aes_core/SB1/n1907 ,
         \U1/aes_core/SB1/n1906 , \U1/aes_core/SB1/n1905 ,
         \U1/aes_core/SB1/n1904 , \U1/aes_core/SB1/n1903 ,
         \U1/aes_core/SB1/n1902 , \U1/aes_core/SB1/n1901 ,
         \U1/aes_core/SB1/n1900 , \U1/aes_core/SB1/n1899 ,
         \U1/aes_core/SB1/n1898 , \U1/aes_core/SB1/n1897 ,
         \U1/aes_core/SB1/n1896 , \U1/aes_core/SB1/n1895 ,
         \U1/aes_core/SB1/n1894 , \U1/aes_core/SB1/n1893 ,
         \U1/aes_core/SB1/n1892 , \U1/aes_core/SB1/n1891 ,
         \U1/aes_core/SB1/n1890 , \U1/aes_core/SB1/n1889 ,
         \U1/aes_core/SB1/n1888 , \U1/aes_core/SB1/n1887 ,
         \U1/aes_core/SB1/n1886 , \U1/aes_core/SB1/n1885 ,
         \U1/aes_core/SB1/n1884 , \U1/aes_core/SB1/n1883 ,
         \U1/aes_core/SB1/n1882 , \U1/aes_core/SB1/n1881 ,
         \U1/aes_core/SB1/n1880 , \U1/aes_core/SB1/n1879 ,
         \U1/aes_core/SB1/n1878 , \U1/aes_core/SB1/n1877 ,
         \U1/aes_core/SB1/n1876 , \U1/aes_core/SB1/n1875 ,
         \U1/aes_core/SB1/n1874 , \U1/aes_core/SB1/n1873 ,
         \U1/aes_core/SB1/n1872 , \U1/aes_core/SB1/n1871 ,
         \U1/aes_core/SB1/n1870 , \U1/aes_core/SB1/n1869 ,
         \U1/aes_core/SB1/n1868 , \U1/aes_core/SB1/n1867 ,
         \U1/aes_core/SB1/n1866 , \U1/aes_core/SB1/n1865 ,
         \U1/aes_core/SB1/n1864 , \U1/aes_core/SB1/n1863 ,
         \U1/aes_core/SB1/n1862 , \U1/aes_core/SB1/n1861 ,
         \U1/aes_core/SB1/n1860 , \U1/aes_core/SB1/n1859 ,
         \U1/aes_core/SB1/n1858 , \U1/aes_core/SB1/n1857 ,
         \U1/aes_core/SB1/n1856 , \U1/aes_core/SB1/n1855 ,
         \U1/aes_core/SB1/n1854 , \U1/aes_core/SB1/n1853 ,
         \U1/aes_core/SB1/n1852 , \U1/aes_core/SB1/n1851 ,
         \U1/aes_core/SB1/n1850 , \U1/aes_core/SB1/n1849 ,
         \U1/aes_core/SB1/n1848 , \U1/aes_core/SB1/n1847 ,
         \U1/aes_core/SB1/n1846 , \U1/aes_core/SB1/n1845 ,
         \U1/aes_core/SB1/n1844 , \U1/aes_core/SB1/n1843 ,
         \U1/aes_core/SB1/n1842 , \U1/aes_core/SB1/n1841 ,
         \U1/aes_core/SB1/n1840 , \U1/aes_core/SB1/n1839 ,
         \U1/aes_core/SB1/n1838 , \U1/aes_core/SB1/n1837 ,
         \U1/aes_core/SB1/n1836 , \U1/aes_core/SB1/n1835 ,
         \U1/aes_core/SB1/n1834 , \U1/aes_core/SB1/n1833 ,
         \U1/aes_core/SB1/n1832 , \U1/aes_core/SB1/n1831 ,
         \U1/aes_core/SB1/n1830 , \U1/aes_core/SB1/n1829 ,
         \U1/aes_core/SB1/n1828 , \U1/aes_core/SB1/n1827 ,
         \U1/aes_core/SB1/n1826 , \U1/aes_core/SB1/n1825 ,
         \U1/aes_core/SB1/n1824 , \U1/aes_core/SB1/n1823 ,
         \U1/aes_core/SB1/n1822 , \U1/aes_core/SB1/n1821 ,
         \U1/aes_core/SB1/n1820 , \U1/aes_core/SB1/n1819 ,
         \U1/aes_core/SB1/n1818 , \U1/aes_core/SB1/n1817 ,
         \U1/aes_core/SB1/n1816 , \U1/aes_core/SB1/n1815 ,
         \U1/aes_core/SB1/n1814 , \U1/aes_core/SB1/n1813 ,
         \U1/aes_core/SB1/n1812 , \U1/aes_core/SB1/n1811 ,
         \U1/aes_core/SB1/n1810 , \U1/aes_core/SB1/n1809 ,
         \U1/aes_core/SB1/n1808 , \U1/aes_core/SB1/n1807 ,
         \U1/aes_core/SB1/n1806 , \U1/aes_core/SB1/n1805 ,
         \U1/aes_core/SB1/n1804 , \U1/aes_core/SB1/n1803 ,
         \U1/aes_core/SB1/n1802 , \U1/aes_core/SB1/n1801 ,
         \U1/aes_core/SB1/n1800 , \U1/aes_core/SB1/n1799 ,
         \U1/aes_core/SB1/n1798 , \U1/aes_core/SB1/n1797 ,
         \U1/aes_core/SB1/n1796 , \U1/aes_core/SB1/n1795 ,
         \U1/aes_core/SB1/n1794 , \U1/aes_core/SB1/n1793 ,
         \U1/aes_core/SB1/n1792 , \U1/aes_core/SB1/n1791 ,
         \U1/aes_core/SB1/n1790 , \U1/aes_core/SB1/n1789 ,
         \U1/aes_core/SB1/n1788 , \U1/aes_core/SB1/n1787 ,
         \U1/aes_core/SB1/n1786 , \U1/aes_core/SB1/n1785 ,
         \U1/aes_core/SB1/n1784 , \U1/aes_core/SB1/n1783 ,
         \U1/aes_core/SB1/n1782 , \U1/aes_core/SB1/n1781 ,
         \U1/aes_core/SB1/n1780 , \U1/aes_core/SB1/n1779 ,
         \U1/aes_core/SB1/n1778 , \U1/aes_core/SB1/n1777 ,
         \U1/aes_core/SB1/n1776 , \U1/aes_core/SB1/n1775 ,
         \U1/aes_core/SB1/n1774 , \U1/aes_core/SB1/n1773 ,
         \U1/aes_core/SB1/n1772 , \U1/aes_core/SB1/n1771 ,
         \U1/aes_core/SB1/n1770 , \U1/aes_core/SB1/n1769 ,
         \U1/aes_core/SB1/n1768 , \U1/aes_core/SB1/n1767 ,
         \U1/aes_core/SB1/n1766 , \U1/aes_core/SB1/n1765 ,
         \U1/aes_core/SB1/n1764 , \U1/aes_core/SB1/n1763 ,
         \U1/aes_core/SB1/n1762 , \U1/aes_core/SB1/n1761 ,
         \U1/aes_core/SB1/n1760 , \U1/aes_core/SB1/n1759 ,
         \U1/aes_core/SB1/n1758 , \U1/aes_core/SB1/n1757 ,
         \U1/aes_core/SB1/n1756 , \U1/aes_core/SB1/n1755 ,
         \U1/aes_core/SB1/n1754 , \U1/aes_core/SB1/n1753 ,
         \U1/aes_core/SB1/n1752 , \U1/aes_core/SB1/n1751 ,
         \U1/aes_core/SB1/n1750 , \U1/aes_core/SB1/n1749 ,
         \U1/aes_core/SB1/n1748 , \U1/aes_core/SB1/n1747 ,
         \U1/aes_core/SB1/n1746 , \U1/aes_core/SB1/n1745 ,
         \U1/aes_core/SB1/n1744 , \U1/aes_core/SB1/n1743 ,
         \U1/aes_core/SB1/n1742 , \U1/aes_core/SB1/n1741 ,
         \U1/aes_core/SB1/n1740 , \U1/aes_core/SB1/n1739 ,
         \U1/aes_core/SB1/n1738 , \U1/aes_core/SB1/n1737 ,
         \U1/aes_core/SB1/n1736 , \U1/aes_core/SB1/n1735 ,
         \U1/aes_core/SB1/n1734 , \U1/aes_core/SB1/n1733 ,
         \U1/aes_core/SB1/n1732 , \U1/aes_core/SB1/n1731 ,
         \U1/aes_core/SB1/n1730 , \U1/aes_core/SB1/n1729 ,
         \U1/aes_core/SB1/n1728 , \U1/aes_core/SB1/n1727 ,
         \U1/aes_core/SB1/n1726 , \U1/aes_core/SB1/n1725 ,
         \U1/aes_core/SB1/n1724 , \U1/aes_core/SB1/n1723 ,
         \U1/aes_core/SB1/n1722 , \U1/aes_core/SB1/n1721 ,
         \U1/aes_core/SB1/n1720 , \U1/aes_core/SB1/n1719 ,
         \U1/aes_core/SB1/n1718 , \U1/aes_core/SB1/n1717 ,
         \U1/aes_core/SB1/n1716 , \U1/aes_core/SB1/n1715 ,
         \U1/aes_core/SB1/n1714 , \U1/aes_core/SB1/n1713 ,
         \U1/aes_core/SB1/n1712 , \U1/aes_core/SB1/n1711 ,
         \U1/aes_core/SB1/n1710 , \U1/aes_core/SB1/n1709 ,
         \U1/aes_core/SB1/n1708 , \U1/aes_core/SB1/n1707 ,
         \U1/aes_core/SB1/n1706 , \U1/aes_core/SB1/n1705 ,
         \U1/aes_core/SB1/n1704 , \U1/aes_core/SB1/n1703 ,
         \U1/aes_core/SB1/n1702 , \U1/aes_core/SB1/n1701 ,
         \U1/aes_core/SB1/n1700 , \U1/aes_core/SB1/n1699 ,
         \U1/aes_core/SB1/n1698 , \U1/aes_core/SB1/n1697 ,
         \U1/aes_core/SB1/n1696 , \U1/aes_core/SB1/n1695 ,
         \U1/aes_core/SB1/n1694 , \U1/aes_core/SB1/n1693 ,
         \U1/aes_core/SB1/n1692 , \U1/aes_core/SB1/n1691 ,
         \U1/aes_core/SB1/n1690 , \U1/aes_core/SB1/n1689 ,
         \U1/aes_core/SB1/n1688 , \U1/aes_core/SB1/n1687 ,
         \U1/aes_core/SB1/n1686 , \U1/aes_core/SB1/n1685 ,
         \U1/aes_core/SB1/n1684 , \U1/aes_core/SB1/n1683 ,
         \U1/aes_core/SB1/n1682 , \U1/aes_core/SB1/n1621 ,
         \U1/aes_core/SB1/n1218 , \U1/aes_core/SB1/n1203 ,
         \U1/aes_core/SB1/n1158 , \U1/aes_core/SB1/n1030 ,
         \U1/aes_core/SB1/n767 , \U1/aes_core/SB1/n752 ,
         \U1/aes_core/SB1/n707 , \U1/aes_core/SB1/n385 ,
         \U1/aes_core/SB2/n3353 , \U1/aes_core/SB2/n3352 ,
         \U1/aes_core/SB2/n3351 , \U1/aes_core/SB2/n3350 ,
         \U1/aes_core/SB2/n3349 , \U1/aes_core/SB2/n3348 ,
         \U1/aes_core/SB2/n3347 , \U1/aes_core/SB2/n3346 ,
         \U1/aes_core/SB2/n3345 , \U1/aes_core/SB2/n3344 ,
         \U1/aes_core/SB2/n3343 , \U1/aes_core/SB2/n3342 ,
         \U1/aes_core/SB2/n3341 , \U1/aes_core/SB2/n3340 ,
         \U1/aes_core/SB2/n3339 , \U1/aes_core/SB2/n3338 ,
         \U1/aes_core/SB2/n3337 , \U1/aes_core/SB2/n3336 ,
         \U1/aes_core/SB2/n3335 , \U1/aes_core/SB2/n3334 ,
         \U1/aes_core/SB2/n3333 , \U1/aes_core/SB2/n3332 ,
         \U1/aes_core/SB2/n3331 , \U1/aes_core/SB2/n3330 ,
         \U1/aes_core/SB2/n3329 , \U1/aes_core/SB2/n3328 ,
         \U1/aes_core/SB2/n3327 , \U1/aes_core/SB2/n3326 ,
         \U1/aes_core/SB2/n3325 , \U1/aes_core/SB2/n3324 ,
         \U1/aes_core/SB2/n3323 , \U1/aes_core/SB2/n3322 ,
         \U1/aes_core/SB2/n3321 , \U1/aes_core/SB2/n3320 ,
         \U1/aes_core/SB2/n3319 , \U1/aes_core/SB2/n3318 ,
         \U1/aes_core/SB2/n3317 , \U1/aes_core/SB2/n3316 ,
         \U1/aes_core/SB2/n3315 , \U1/aes_core/SB2/n3314 ,
         \U1/aes_core/SB2/n3313 , \U1/aes_core/SB2/n3312 ,
         \U1/aes_core/SB2/n3311 , \U1/aes_core/SB2/n3310 ,
         \U1/aes_core/SB2/n3309 , \U1/aes_core/SB2/n3308 ,
         \U1/aes_core/SB2/n3307 , \U1/aes_core/SB2/n3306 ,
         \U1/aes_core/SB2/n3305 , \U1/aes_core/SB2/n3304 ,
         \U1/aes_core/SB2/n3303 , \U1/aes_core/SB2/n3302 ,
         \U1/aes_core/SB2/n3301 , \U1/aes_core/SB2/n3300 ,
         \U1/aes_core/SB2/n3299 , \U1/aes_core/SB2/n3298 ,
         \U1/aes_core/SB2/n3297 , \U1/aes_core/SB2/n3296 ,
         \U1/aes_core/SB2/n3295 , \U1/aes_core/SB2/n3294 ,
         \U1/aes_core/SB2/n3293 , \U1/aes_core/SB2/n3292 ,
         \U1/aes_core/SB2/n3291 , \U1/aes_core/SB2/n3290 ,
         \U1/aes_core/SB2/n3289 , \U1/aes_core/SB2/n3288 ,
         \U1/aes_core/SB2/n3287 , \U1/aes_core/SB2/n3286 ,
         \U1/aes_core/SB2/n3285 , \U1/aes_core/SB2/n3284 ,
         \U1/aes_core/SB2/n3283 , \U1/aes_core/SB2/n3282 ,
         \U1/aes_core/SB2/n3281 , \U1/aes_core/SB2/n3280 ,
         \U1/aes_core/SB2/n3279 , \U1/aes_core/SB2/n3278 ,
         \U1/aes_core/SB2/n3277 , \U1/aes_core/SB2/n3276 ,
         \U1/aes_core/SB2/n3275 , \U1/aes_core/SB2/n3274 ,
         \U1/aes_core/SB2/n3273 , \U1/aes_core/SB2/n3272 ,
         \U1/aes_core/SB2/n3271 , \U1/aes_core/SB2/n3270 ,
         \U1/aes_core/SB2/n3269 , \U1/aes_core/SB2/n3268 ,
         \U1/aes_core/SB2/n3267 , \U1/aes_core/SB2/n3266 ,
         \U1/aes_core/SB2/n3265 , \U1/aes_core/SB2/n3264 ,
         \U1/aes_core/SB2/n3263 , \U1/aes_core/SB2/n3262 ,
         \U1/aes_core/SB2/n3261 , \U1/aes_core/SB2/n3260 ,
         \U1/aes_core/SB2/n3259 , \U1/aes_core/SB2/n3258 ,
         \U1/aes_core/SB2/n3257 , \U1/aes_core/SB2/n3256 ,
         \U1/aes_core/SB2/n3255 , \U1/aes_core/SB2/n3254 ,
         \U1/aes_core/SB2/n3253 , \U1/aes_core/SB2/n3252 ,
         \U1/aes_core/SB2/n3251 , \U1/aes_core/SB2/n3250 ,
         \U1/aes_core/SB2/n3249 , \U1/aes_core/SB2/n3248 ,
         \U1/aes_core/SB2/n3247 , \U1/aes_core/SB2/n3246 ,
         \U1/aes_core/SB2/n3245 , \U1/aes_core/SB2/n3244 ,
         \U1/aes_core/SB2/n3243 , \U1/aes_core/SB2/n3242 ,
         \U1/aes_core/SB2/n3241 , \U1/aes_core/SB2/n3240 ,
         \U1/aes_core/SB2/n3239 , \U1/aes_core/SB2/n3238 ,
         \U1/aes_core/SB2/n3237 , \U1/aes_core/SB2/n3236 ,
         \U1/aes_core/SB2/n3235 , \U1/aes_core/SB2/n3234 ,
         \U1/aes_core/SB2/n3233 , \U1/aes_core/SB2/n3232 ,
         \U1/aes_core/SB2/n3231 , \U1/aes_core/SB2/n3230 ,
         \U1/aes_core/SB2/n3229 , \U1/aes_core/SB2/n3228 ,
         \U1/aes_core/SB2/n3227 , \U1/aes_core/SB2/n3226 ,
         \U1/aes_core/SB2/n3225 , \U1/aes_core/SB2/n3224 ,
         \U1/aes_core/SB2/n3223 , \U1/aes_core/SB2/n3222 ,
         \U1/aes_core/SB2/n3221 , \U1/aes_core/SB2/n3220 ,
         \U1/aes_core/SB2/n3219 , \U1/aes_core/SB2/n3218 ,
         \U1/aes_core/SB2/n3217 , \U1/aes_core/SB2/n3216 ,
         \U1/aes_core/SB2/n3215 , \U1/aes_core/SB2/n3214 ,
         \U1/aes_core/SB2/n3213 , \U1/aes_core/SB2/n3212 ,
         \U1/aes_core/SB2/n3211 , \U1/aes_core/SB2/n3210 ,
         \U1/aes_core/SB2/n3209 , \U1/aes_core/SB2/n3208 ,
         \U1/aes_core/SB2/n3207 , \U1/aes_core/SB2/n3206 ,
         \U1/aes_core/SB2/n3205 , \U1/aes_core/SB2/n3204 ,
         \U1/aes_core/SB2/n3203 , \U1/aes_core/SB2/n3202 ,
         \U1/aes_core/SB2/n3201 , \U1/aes_core/SB2/n3200 ,
         \U1/aes_core/SB2/n3199 , \U1/aes_core/SB2/n3198 ,
         \U1/aes_core/SB2/n3197 , \U1/aes_core/SB2/n3196 ,
         \U1/aes_core/SB2/n3195 , \U1/aes_core/SB2/n3194 ,
         \U1/aes_core/SB2/n3193 , \U1/aes_core/SB2/n3192 ,
         \U1/aes_core/SB2/n3191 , \U1/aes_core/SB2/n3190 ,
         \U1/aes_core/SB2/n3189 , \U1/aes_core/SB2/n3188 ,
         \U1/aes_core/SB2/n3187 , \U1/aes_core/SB2/n3186 ,
         \U1/aes_core/SB2/n3185 , \U1/aes_core/SB2/n3184 ,
         \U1/aes_core/SB2/n3183 , \U1/aes_core/SB2/n3182 ,
         \U1/aes_core/SB2/n3181 , \U1/aes_core/SB2/n3180 ,
         \U1/aes_core/SB2/n3179 , \U1/aes_core/SB2/n3178 ,
         \U1/aes_core/SB2/n3177 , \U1/aes_core/SB2/n3176 ,
         \U1/aes_core/SB2/n3175 , \U1/aes_core/SB2/n3174 ,
         \U1/aes_core/SB2/n3173 , \U1/aes_core/SB2/n3172 ,
         \U1/aes_core/SB2/n3171 , \U1/aes_core/SB2/n3170 ,
         \U1/aes_core/SB2/n3169 , \U1/aes_core/SB2/n3168 ,
         \U1/aes_core/SB2/n3167 , \U1/aes_core/SB2/n3166 ,
         \U1/aes_core/SB2/n3165 , \U1/aes_core/SB2/n3164 ,
         \U1/aes_core/SB2/n3163 , \U1/aes_core/SB2/n3162 ,
         \U1/aes_core/SB2/n3161 , \U1/aes_core/SB2/n3160 ,
         \U1/aes_core/SB2/n3159 , \U1/aes_core/SB2/n3158 ,
         \U1/aes_core/SB2/n3157 , \U1/aes_core/SB2/n3156 ,
         \U1/aes_core/SB2/n3155 , \U1/aes_core/SB2/n3154 ,
         \U1/aes_core/SB2/n3153 , \U1/aes_core/SB2/n3152 ,
         \U1/aes_core/SB2/n3151 , \U1/aes_core/SB2/n3150 ,
         \U1/aes_core/SB2/n3149 , \U1/aes_core/SB2/n3148 ,
         \U1/aes_core/SB2/n3147 , \U1/aes_core/SB2/n3146 ,
         \U1/aes_core/SB2/n3145 , \U1/aes_core/SB2/n3144 ,
         \U1/aes_core/SB2/n3143 , \U1/aes_core/SB2/n3142 ,
         \U1/aes_core/SB2/n3141 , \U1/aes_core/SB2/n3140 ,
         \U1/aes_core/SB2/n3139 , \U1/aes_core/SB2/n3138 ,
         \U1/aes_core/SB2/n3137 , \U1/aes_core/SB2/n3136 ,
         \U1/aes_core/SB2/n3135 , \U1/aes_core/SB2/n3134 ,
         \U1/aes_core/SB2/n3133 , \U1/aes_core/SB2/n3132 ,
         \U1/aes_core/SB2/n3131 , \U1/aes_core/SB2/n3130 ,
         \U1/aes_core/SB2/n3129 , \U1/aes_core/SB2/n3128 ,
         \U1/aes_core/SB2/n3127 , \U1/aes_core/SB2/n3126 ,
         \U1/aes_core/SB2/n3125 , \U1/aes_core/SB2/n3124 ,
         \U1/aes_core/SB2/n3123 , \U1/aes_core/SB2/n3122 ,
         \U1/aes_core/SB2/n3121 , \U1/aes_core/SB2/n3120 ,
         \U1/aes_core/SB2/n3119 , \U1/aes_core/SB2/n3118 ,
         \U1/aes_core/SB2/n3117 , \U1/aes_core/SB2/n3116 ,
         \U1/aes_core/SB2/n3115 , \U1/aes_core/SB2/n3114 ,
         \U1/aes_core/SB2/n3113 , \U1/aes_core/SB2/n3112 ,
         \U1/aes_core/SB2/n3111 , \U1/aes_core/SB2/n3110 ,
         \U1/aes_core/SB2/n3109 , \U1/aes_core/SB2/n3108 ,
         \U1/aes_core/SB2/n3107 , \U1/aes_core/SB2/n3106 ,
         \U1/aes_core/SB2/n3105 , \U1/aes_core/SB2/n3104 ,
         \U1/aes_core/SB2/n3103 , \U1/aes_core/SB2/n3102 ,
         \U1/aes_core/SB2/n3101 , \U1/aes_core/SB2/n3100 ,
         \U1/aes_core/SB2/n3099 , \U1/aes_core/SB2/n3098 ,
         \U1/aes_core/SB2/n3097 , \U1/aes_core/SB2/n3096 ,
         \U1/aes_core/SB2/n3095 , \U1/aes_core/SB2/n3094 ,
         \U1/aes_core/SB2/n3093 , \U1/aes_core/SB2/n3092 ,
         \U1/aes_core/SB2/n3091 , \U1/aes_core/SB2/n3090 ,
         \U1/aes_core/SB2/n3089 , \U1/aes_core/SB2/n3088 ,
         \U1/aes_core/SB2/n3087 , \U1/aes_core/SB2/n3086 ,
         \U1/aes_core/SB2/n3085 , \U1/aes_core/SB2/n3084 ,
         \U1/aes_core/SB2/n3083 , \U1/aes_core/SB2/n3082 ,
         \U1/aes_core/SB2/n3081 , \U1/aes_core/SB2/n3080 ,
         \U1/aes_core/SB2/n3079 , \U1/aes_core/SB2/n3078 ,
         \U1/aes_core/SB2/n3077 , \U1/aes_core/SB2/n3076 ,
         \U1/aes_core/SB2/n3075 , \U1/aes_core/SB2/n3074 ,
         \U1/aes_core/SB2/n3073 , \U1/aes_core/SB2/n3072 ,
         \U1/aes_core/SB2/n3071 , \U1/aes_core/SB2/n3070 ,
         \U1/aes_core/SB2/n3069 , \U1/aes_core/SB2/n3068 ,
         \U1/aes_core/SB2/n3067 , \U1/aes_core/SB2/n3066 ,
         \U1/aes_core/SB2/n3065 , \U1/aes_core/SB2/n3064 ,
         \U1/aes_core/SB2/n3063 , \U1/aes_core/SB2/n3062 ,
         \U1/aes_core/SB2/n3061 , \U1/aes_core/SB2/n3060 ,
         \U1/aes_core/SB2/n3059 , \U1/aes_core/SB2/n3058 ,
         \U1/aes_core/SB2/n3057 , \U1/aes_core/SB2/n3056 ,
         \U1/aes_core/SB2/n3055 , \U1/aes_core/SB2/n3054 ,
         \U1/aes_core/SB2/n3053 , \U1/aes_core/SB2/n3052 ,
         \U1/aes_core/SB2/n3051 , \U1/aes_core/SB2/n3050 ,
         \U1/aes_core/SB2/n3049 , \U1/aes_core/SB2/n3048 ,
         \U1/aes_core/SB2/n3047 , \U1/aes_core/SB2/n3046 ,
         \U1/aes_core/SB2/n3045 , \U1/aes_core/SB2/n3044 ,
         \U1/aes_core/SB2/n3043 , \U1/aes_core/SB2/n3042 ,
         \U1/aes_core/SB2/n3041 , \U1/aes_core/SB2/n3040 ,
         \U1/aes_core/SB2/n3039 , \U1/aes_core/SB2/n3038 ,
         \U1/aes_core/SB2/n3037 , \U1/aes_core/SB2/n3036 ,
         \U1/aes_core/SB2/n3035 , \U1/aes_core/SB2/n3034 ,
         \U1/aes_core/SB2/n3033 , \U1/aes_core/SB2/n3032 ,
         \U1/aes_core/SB2/n3031 , \U1/aes_core/SB2/n3030 ,
         \U1/aes_core/SB2/n3029 , \U1/aes_core/SB2/n3028 ,
         \U1/aes_core/SB2/n3027 , \U1/aes_core/SB2/n3026 ,
         \U1/aes_core/SB2/n3025 , \U1/aes_core/SB2/n3024 ,
         \U1/aes_core/SB2/n3023 , \U1/aes_core/SB2/n3022 ,
         \U1/aes_core/SB2/n3021 , \U1/aes_core/SB2/n3020 ,
         \U1/aes_core/SB2/n3019 , \U1/aes_core/SB2/n3018 ,
         \U1/aes_core/SB2/n3017 , \U1/aes_core/SB2/n3016 ,
         \U1/aes_core/SB2/n3015 , \U1/aes_core/SB2/n3014 ,
         \U1/aes_core/SB2/n3013 , \U1/aes_core/SB2/n3012 ,
         \U1/aes_core/SB2/n3011 , \U1/aes_core/SB2/n3010 ,
         \U1/aes_core/SB2/n3009 , \U1/aes_core/SB2/n3008 ,
         \U1/aes_core/SB2/n3007 , \U1/aes_core/SB2/n3006 ,
         \U1/aes_core/SB2/n3005 , \U1/aes_core/SB2/n3004 ,
         \U1/aes_core/SB2/n3003 , \U1/aes_core/SB2/n3002 ,
         \U1/aes_core/SB2/n3001 , \U1/aes_core/SB2/n3000 ,
         \U1/aes_core/SB2/n2999 , \U1/aes_core/SB2/n2998 ,
         \U1/aes_core/SB2/n2997 , \U1/aes_core/SB2/n2996 ,
         \U1/aes_core/SB2/n2995 , \U1/aes_core/SB2/n2994 ,
         \U1/aes_core/SB2/n2993 , \U1/aes_core/SB2/n2992 ,
         \U1/aes_core/SB2/n2991 , \U1/aes_core/SB2/n2990 ,
         \U1/aes_core/SB2/n2989 , \U1/aes_core/SB2/n2988 ,
         \U1/aes_core/SB2/n2987 , \U1/aes_core/SB2/n2986 ,
         \U1/aes_core/SB2/n2985 , \U1/aes_core/SB2/n2984 ,
         \U1/aes_core/SB2/n2983 , \U1/aes_core/SB2/n2982 ,
         \U1/aes_core/SB2/n2981 , \U1/aes_core/SB2/n2980 ,
         \U1/aes_core/SB2/n2979 , \U1/aes_core/SB2/n2978 ,
         \U1/aes_core/SB2/n2977 , \U1/aes_core/SB2/n2976 ,
         \U1/aes_core/SB2/n2975 , \U1/aes_core/SB2/n2974 ,
         \U1/aes_core/SB2/n2973 , \U1/aes_core/SB2/n2972 ,
         \U1/aes_core/SB2/n2971 , \U1/aes_core/SB2/n2970 ,
         \U1/aes_core/SB2/n2969 , \U1/aes_core/SB2/n2968 ,
         \U1/aes_core/SB2/n2967 , \U1/aes_core/SB2/n2966 ,
         \U1/aes_core/SB2/n2965 , \U1/aes_core/SB2/n2964 ,
         \U1/aes_core/SB2/n2963 , \U1/aes_core/SB2/n2962 ,
         \U1/aes_core/SB2/n2961 , \U1/aes_core/SB2/n2960 ,
         \U1/aes_core/SB2/n2959 , \U1/aes_core/SB2/n2958 ,
         \U1/aes_core/SB2/n2957 , \U1/aes_core/SB2/n2956 ,
         \U1/aes_core/SB2/n2955 , \U1/aes_core/SB2/n2954 ,
         \U1/aes_core/SB2/n2953 , \U1/aes_core/SB2/n2952 ,
         \U1/aes_core/SB2/n2951 , \U1/aes_core/SB2/n2950 ,
         \U1/aes_core/SB2/n2949 , \U1/aes_core/SB2/n2948 ,
         \U1/aes_core/SB2/n2947 , \U1/aes_core/SB2/n2946 ,
         \U1/aes_core/SB2/n2945 , \U1/aes_core/SB2/n2944 ,
         \U1/aes_core/SB2/n2943 , \U1/aes_core/SB2/n2942 ,
         \U1/aes_core/SB2/n2941 , \U1/aes_core/SB2/n2940 ,
         \U1/aes_core/SB2/n2939 , \U1/aes_core/SB2/n2938 ,
         \U1/aes_core/SB2/n2937 , \U1/aes_core/SB2/n2936 ,
         \U1/aes_core/SB2/n2935 , \U1/aes_core/SB2/n2934 ,
         \U1/aes_core/SB2/n2933 , \U1/aes_core/SB2/n2932 ,
         \U1/aes_core/SB2/n2931 , \U1/aes_core/SB2/n2930 ,
         \U1/aes_core/SB2/n2929 , \U1/aes_core/SB2/n2928 ,
         \U1/aes_core/SB2/n2927 , \U1/aes_core/SB2/n2926 ,
         \U1/aes_core/SB2/n2925 , \U1/aes_core/SB2/n2924 ,
         \U1/aes_core/SB2/n2923 , \U1/aes_core/SB2/n2922 ,
         \U1/aes_core/SB2/n2921 , \U1/aes_core/SB2/n2920 ,
         \U1/aes_core/SB2/n2919 , \U1/aes_core/SB2/n2918 ,
         \U1/aes_core/SB2/n2917 , \U1/aes_core/SB2/n2916 ,
         \U1/aes_core/SB2/n2915 , \U1/aes_core/SB2/n2914 ,
         \U1/aes_core/SB2/n2913 , \U1/aes_core/SB2/n2912 ,
         \U1/aes_core/SB2/n2911 , \U1/aes_core/SB2/n2910 ,
         \U1/aes_core/SB2/n2909 , \U1/aes_core/SB2/n2908 ,
         \U1/aes_core/SB2/n2907 , \U1/aes_core/SB2/n2906 ,
         \U1/aes_core/SB2/n2905 , \U1/aes_core/SB2/n2904 ,
         \U1/aes_core/SB2/n2903 , \U1/aes_core/SB2/n2902 ,
         \U1/aes_core/SB2/n2901 , \U1/aes_core/SB2/n2900 ,
         \U1/aes_core/SB2/n2899 , \U1/aes_core/SB2/n2898 ,
         \U1/aes_core/SB2/n2897 , \U1/aes_core/SB2/n2896 ,
         \U1/aes_core/SB2/n2895 , \U1/aes_core/SB2/n2894 ,
         \U1/aes_core/SB2/n2893 , \U1/aes_core/SB2/n2892 ,
         \U1/aes_core/SB2/n2891 , \U1/aes_core/SB2/n2890 ,
         \U1/aes_core/SB2/n2889 , \U1/aes_core/SB2/n2888 ,
         \U1/aes_core/SB2/n2887 , \U1/aes_core/SB2/n2886 ,
         \U1/aes_core/SB2/n2885 , \U1/aes_core/SB2/n2884 ,
         \U1/aes_core/SB2/n2883 , \U1/aes_core/SB2/n2882 ,
         \U1/aes_core/SB2/n2881 , \U1/aes_core/SB2/n2880 ,
         \U1/aes_core/SB2/n2879 , \U1/aes_core/SB2/n2878 ,
         \U1/aes_core/SB2/n2877 , \U1/aes_core/SB2/n2876 ,
         \U1/aes_core/SB2/n2875 , \U1/aes_core/SB2/n2874 ,
         \U1/aes_core/SB2/n2873 , \U1/aes_core/SB2/n2872 ,
         \U1/aes_core/SB2/n2871 , \U1/aes_core/SB2/n2870 ,
         \U1/aes_core/SB2/n2869 , \U1/aes_core/SB2/n2868 ,
         \U1/aes_core/SB2/n2867 , \U1/aes_core/SB2/n2866 ,
         \U1/aes_core/SB2/n2865 , \U1/aes_core/SB2/n2864 ,
         \U1/aes_core/SB2/n2863 , \U1/aes_core/SB2/n2862 ,
         \U1/aes_core/SB2/n2861 , \U1/aes_core/SB2/n2860 ,
         \U1/aes_core/SB2/n2859 , \U1/aes_core/SB2/n2858 ,
         \U1/aes_core/SB2/n2857 , \U1/aes_core/SB2/n2856 ,
         \U1/aes_core/SB2/n2855 , \U1/aes_core/SB2/n2854 ,
         \U1/aes_core/SB2/n2853 , \U1/aes_core/SB2/n2852 ,
         \U1/aes_core/SB2/n2851 , \U1/aes_core/SB2/n2850 ,
         \U1/aes_core/SB2/n2849 , \U1/aes_core/SB2/n2848 ,
         \U1/aes_core/SB2/n2847 , \U1/aes_core/SB2/n2846 ,
         \U1/aes_core/SB2/n2845 , \U1/aes_core/SB2/n2844 ,
         \U1/aes_core/SB2/n2843 , \U1/aes_core/SB2/n2842 ,
         \U1/aes_core/SB2/n2841 , \U1/aes_core/SB2/n2840 ,
         \U1/aes_core/SB2/n2839 , \U1/aes_core/SB2/n2838 ,
         \U1/aes_core/SB2/n2837 , \U1/aes_core/SB2/n2836 ,
         \U1/aes_core/SB2/n2835 , \U1/aes_core/SB2/n2834 ,
         \U1/aes_core/SB2/n2833 , \U1/aes_core/SB2/n2832 ,
         \U1/aes_core/SB2/n2831 , \U1/aes_core/SB2/n2830 ,
         \U1/aes_core/SB2/n2829 , \U1/aes_core/SB2/n2828 ,
         \U1/aes_core/SB2/n2827 , \U1/aes_core/SB2/n2826 ,
         \U1/aes_core/SB2/n2825 , \U1/aes_core/SB2/n2824 ,
         \U1/aes_core/SB2/n2823 , \U1/aes_core/SB2/n2822 ,
         \U1/aes_core/SB2/n2821 , \U1/aes_core/SB2/n2820 ,
         \U1/aes_core/SB2/n2819 , \U1/aes_core/SB2/n2818 ,
         \U1/aes_core/SB2/n2817 , \U1/aes_core/SB2/n2816 ,
         \U1/aes_core/SB2/n2815 , \U1/aes_core/SB2/n2814 ,
         \U1/aes_core/SB2/n2813 , \U1/aes_core/SB2/n2812 ,
         \U1/aes_core/SB2/n2811 , \U1/aes_core/SB2/n2810 ,
         \U1/aes_core/SB2/n2809 , \U1/aes_core/SB2/n2808 ,
         \U1/aes_core/SB2/n2807 , \U1/aes_core/SB2/n2806 ,
         \U1/aes_core/SB2/n2805 , \U1/aes_core/SB2/n2804 ,
         \U1/aes_core/SB2/n2803 , \U1/aes_core/SB2/n2802 ,
         \U1/aes_core/SB2/n2801 , \U1/aes_core/SB2/n2800 ,
         \U1/aes_core/SB2/n2799 , \U1/aes_core/SB2/n2798 ,
         \U1/aes_core/SB2/n2797 , \U1/aes_core/SB2/n2796 ,
         \U1/aes_core/SB2/n2795 , \U1/aes_core/SB2/n2794 ,
         \U1/aes_core/SB2/n2793 , \U1/aes_core/SB2/n2792 ,
         \U1/aes_core/SB2/n2791 , \U1/aes_core/SB2/n2790 ,
         \U1/aes_core/SB2/n2789 , \U1/aes_core/SB2/n2788 ,
         \U1/aes_core/SB2/n2787 , \U1/aes_core/SB2/n2786 ,
         \U1/aes_core/SB2/n2785 , \U1/aes_core/SB2/n2784 ,
         \U1/aes_core/SB2/n2783 , \U1/aes_core/SB2/n2782 ,
         \U1/aes_core/SB2/n2781 , \U1/aes_core/SB2/n2780 ,
         \U1/aes_core/SB2/n2779 , \U1/aes_core/SB2/n2778 ,
         \U1/aes_core/SB2/n2777 , \U1/aes_core/SB2/n2776 ,
         \U1/aes_core/SB2/n2775 , \U1/aes_core/SB2/n2774 ,
         \U1/aes_core/SB2/n2773 , \U1/aes_core/SB2/n2772 ,
         \U1/aes_core/SB2/n2771 , \U1/aes_core/SB2/n2770 ,
         \U1/aes_core/SB2/n2769 , \U1/aes_core/SB2/n2768 ,
         \U1/aes_core/SB2/n2767 , \U1/aes_core/SB2/n2766 ,
         \U1/aes_core/SB2/n2765 , \U1/aes_core/SB2/n2764 ,
         \U1/aes_core/SB2/n2763 , \U1/aes_core/SB2/n2762 ,
         \U1/aes_core/SB2/n2761 , \U1/aes_core/SB2/n2760 ,
         \U1/aes_core/SB2/n2759 , \U1/aes_core/SB2/n2758 ,
         \U1/aes_core/SB2/n2757 , \U1/aes_core/SB2/n2756 ,
         \U1/aes_core/SB2/n2755 , \U1/aes_core/SB2/n2754 ,
         \U1/aes_core/SB2/n2753 , \U1/aes_core/SB2/n2752 ,
         \U1/aes_core/SB2/n2751 , \U1/aes_core/SB2/n2750 ,
         \U1/aes_core/SB2/n2749 , \U1/aes_core/SB2/n2748 ,
         \U1/aes_core/SB2/n2747 , \U1/aes_core/SB2/n2746 ,
         \U1/aes_core/SB2/n2745 , \U1/aes_core/SB2/n2744 ,
         \U1/aes_core/SB2/n2743 , \U1/aes_core/SB2/n2742 ,
         \U1/aes_core/SB2/n2741 , \U1/aes_core/SB2/n2740 ,
         \U1/aes_core/SB2/n2739 , \U1/aes_core/SB2/n2738 ,
         \U1/aes_core/SB2/n2737 , \U1/aes_core/SB2/n2736 ,
         \U1/aes_core/SB2/n2735 , \U1/aes_core/SB2/n2734 ,
         \U1/aes_core/SB2/n2733 , \U1/aes_core/SB2/n2732 ,
         \U1/aes_core/SB2/n2731 , \U1/aes_core/SB2/n2730 ,
         \U1/aes_core/SB2/n2729 , \U1/aes_core/SB2/n2728 ,
         \U1/aes_core/SB2/n2727 , \U1/aes_core/SB2/n2726 ,
         \U1/aes_core/SB2/n2725 , \U1/aes_core/SB2/n2724 ,
         \U1/aes_core/SB2/n2723 , \U1/aes_core/SB2/n2722 ,
         \U1/aes_core/SB2/n2721 , \U1/aes_core/SB2/n2720 ,
         \U1/aes_core/SB2/n2719 , \U1/aes_core/SB2/n2718 ,
         \U1/aes_core/SB2/n2717 , \U1/aes_core/SB2/n2716 ,
         \U1/aes_core/SB2/n2715 , \U1/aes_core/SB2/n2714 ,
         \U1/aes_core/SB2/n2713 , \U1/aes_core/SB2/n2712 ,
         \U1/aes_core/SB2/n2711 , \U1/aes_core/SB2/n2710 ,
         \U1/aes_core/SB2/n2709 , \U1/aes_core/SB2/n2708 ,
         \U1/aes_core/SB2/n2707 , \U1/aes_core/SB2/n2706 ,
         \U1/aes_core/SB2/n2705 , \U1/aes_core/SB2/n2704 ,
         \U1/aes_core/SB2/n2703 , \U1/aes_core/SB2/n2702 ,
         \U1/aes_core/SB2/n2701 , \U1/aes_core/SB2/n2700 ,
         \U1/aes_core/SB2/n2699 , \U1/aes_core/SB2/n2698 ,
         \U1/aes_core/SB2/n2697 , \U1/aes_core/SB2/n2696 ,
         \U1/aes_core/SB2/n2695 , \U1/aes_core/SB2/n2694 ,
         \U1/aes_core/SB2/n2693 , \U1/aes_core/SB2/n2692 ,
         \U1/aes_core/SB2/n2691 , \U1/aes_core/SB2/n2690 ,
         \U1/aes_core/SB2/n2689 , \U1/aes_core/SB2/n2688 ,
         \U1/aes_core/SB2/n2687 , \U1/aes_core/SB2/n2686 ,
         \U1/aes_core/SB2/n2685 , \U1/aes_core/SB2/n2684 ,
         \U1/aes_core/SB2/n2683 , \U1/aes_core/SB2/n2682 ,
         \U1/aes_core/SB2/n2681 , \U1/aes_core/SB2/n2680 ,
         \U1/aes_core/SB2/n2679 , \U1/aes_core/SB2/n2678 ,
         \U1/aes_core/SB2/n2677 , \U1/aes_core/SB2/n2676 ,
         \U1/aes_core/SB2/n2675 , \U1/aes_core/SB2/n2674 ,
         \U1/aes_core/SB2/n2673 , \U1/aes_core/SB2/n2672 ,
         \U1/aes_core/SB2/n2671 , \U1/aes_core/SB2/n2670 ,
         \U1/aes_core/SB2/n2669 , \U1/aes_core/SB2/n2668 ,
         \U1/aes_core/SB2/n2667 , \U1/aes_core/SB2/n2666 ,
         \U1/aes_core/SB2/n2665 , \U1/aes_core/SB2/n2664 ,
         \U1/aes_core/SB2/n2663 , \U1/aes_core/SB2/n2662 ,
         \U1/aes_core/SB2/n2661 , \U1/aes_core/SB2/n2660 ,
         \U1/aes_core/SB2/n2659 , \U1/aes_core/SB2/n2658 ,
         \U1/aes_core/SB2/n2657 , \U1/aes_core/SB2/n2656 ,
         \U1/aes_core/SB2/n2655 , \U1/aes_core/SB2/n2654 ,
         \U1/aes_core/SB2/n2653 , \U1/aes_core/SB2/n2652 ,
         \U1/aes_core/SB2/n2651 , \U1/aes_core/SB2/n2650 ,
         \U1/aes_core/SB2/n2649 , \U1/aes_core/SB2/n2648 ,
         \U1/aes_core/SB2/n2647 , \U1/aes_core/SB2/n2646 ,
         \U1/aes_core/SB2/n2645 , \U1/aes_core/SB2/n2644 ,
         \U1/aes_core/SB2/n2643 , \U1/aes_core/SB2/n2642 ,
         \U1/aes_core/SB2/n2641 , \U1/aes_core/SB2/n2640 ,
         \U1/aes_core/SB2/n2639 , \U1/aes_core/SB2/n2638 ,
         \U1/aes_core/SB2/n2637 , \U1/aes_core/SB2/n2636 ,
         \U1/aes_core/SB2/n2635 , \U1/aes_core/SB2/n2634 ,
         \U1/aes_core/SB2/n2633 , \U1/aes_core/SB2/n2632 ,
         \U1/aes_core/SB2/n2631 , \U1/aes_core/SB2/n2630 ,
         \U1/aes_core/SB2/n2629 , \U1/aes_core/SB2/n2628 ,
         \U1/aes_core/SB2/n2627 , \U1/aes_core/SB2/n2626 ,
         \U1/aes_core/SB2/n2625 , \U1/aes_core/SB2/n2624 ,
         \U1/aes_core/SB2/n2623 , \U1/aes_core/SB2/n2622 ,
         \U1/aes_core/SB2/n2621 , \U1/aes_core/SB2/n2620 ,
         \U1/aes_core/SB2/n2619 , \U1/aes_core/SB2/n2618 ,
         \U1/aes_core/SB2/n2617 , \U1/aes_core/SB2/n2616 ,
         \U1/aes_core/SB2/n2615 , \U1/aes_core/SB2/n2614 ,
         \U1/aes_core/SB2/n2613 , \U1/aes_core/SB2/n2612 ,
         \U1/aes_core/SB2/n2611 , \U1/aes_core/SB2/n2610 ,
         \U1/aes_core/SB2/n2609 , \U1/aes_core/SB2/n2608 ,
         \U1/aes_core/SB2/n2607 , \U1/aes_core/SB2/n2606 ,
         \U1/aes_core/SB2/n2605 , \U1/aes_core/SB2/n2604 ,
         \U1/aes_core/SB2/n2603 , \U1/aes_core/SB2/n2602 ,
         \U1/aes_core/SB2/n2601 , \U1/aes_core/SB2/n2600 ,
         \U1/aes_core/SB2/n2599 , \U1/aes_core/SB2/n2598 ,
         \U1/aes_core/SB2/n2597 , \U1/aes_core/SB2/n2596 ,
         \U1/aes_core/SB2/n2595 , \U1/aes_core/SB2/n2594 ,
         \U1/aes_core/SB2/n2593 , \U1/aes_core/SB2/n2592 ,
         \U1/aes_core/SB2/n2591 , \U1/aes_core/SB2/n2590 ,
         \U1/aes_core/SB2/n2589 , \U1/aes_core/SB2/n2588 ,
         \U1/aes_core/SB2/n2587 , \U1/aes_core/SB2/n2586 ,
         \U1/aes_core/SB2/n2585 , \U1/aes_core/SB2/n2584 ,
         \U1/aes_core/SB2/n2583 , \U1/aes_core/SB2/n2582 ,
         \U1/aes_core/SB2/n2581 , \U1/aes_core/SB2/n2580 ,
         \U1/aes_core/SB2/n2579 , \U1/aes_core/SB2/n2578 ,
         \U1/aes_core/SB2/n2577 , \U1/aes_core/SB2/n2576 ,
         \U1/aes_core/SB2/n2575 , \U1/aes_core/SB2/n2574 ,
         \U1/aes_core/SB2/n2573 , \U1/aes_core/SB2/n2572 ,
         \U1/aes_core/SB2/n2571 , \U1/aes_core/SB2/n2570 ,
         \U1/aes_core/SB2/n2569 , \U1/aes_core/SB2/n2568 ,
         \U1/aes_core/SB2/n2567 , \U1/aes_core/SB2/n2566 ,
         \U1/aes_core/SB2/n2565 , \U1/aes_core/SB2/n2564 ,
         \U1/aes_core/SB2/n2563 , \U1/aes_core/SB2/n2562 ,
         \U1/aes_core/SB2/n2561 , \U1/aes_core/SB2/n2560 ,
         \U1/aes_core/SB2/n2559 , \U1/aes_core/SB2/n2558 ,
         \U1/aes_core/SB2/n2557 , \U1/aes_core/SB2/n2556 ,
         \U1/aes_core/SB2/n2555 , \U1/aes_core/SB2/n2554 ,
         \U1/aes_core/SB2/n2553 , \U1/aes_core/SB2/n2552 ,
         \U1/aes_core/SB2/n2551 , \U1/aes_core/SB2/n2550 ,
         \U1/aes_core/SB2/n2549 , \U1/aes_core/SB2/n2548 ,
         \U1/aes_core/SB2/n2547 , \U1/aes_core/SB2/n2546 ,
         \U1/aes_core/SB2/n2545 , \U1/aes_core/SB2/n2544 ,
         \U1/aes_core/SB2/n2543 , \U1/aes_core/SB2/n2542 ,
         \U1/aes_core/SB2/n2541 , \U1/aes_core/SB2/n2540 ,
         \U1/aes_core/SB2/n2539 , \U1/aes_core/SB2/n2538 ,
         \U1/aes_core/SB2/n2537 , \U1/aes_core/SB2/n2536 ,
         \U1/aes_core/SB2/n2535 , \U1/aes_core/SB2/n2534 ,
         \U1/aes_core/SB2/n2533 , \U1/aes_core/SB2/n2532 ,
         \U1/aes_core/SB2/n2531 , \U1/aes_core/SB2/n2530 ,
         \U1/aes_core/SB2/n2529 , \U1/aes_core/SB2/n2528 ,
         \U1/aes_core/SB2/n2527 , \U1/aes_core/SB2/n2526 ,
         \U1/aes_core/SB2/n2525 , \U1/aes_core/SB2/n2524 ,
         \U1/aes_core/SB2/n2523 , \U1/aes_core/SB2/n2522 ,
         \U1/aes_core/SB2/n2521 , \U1/aes_core/SB2/n2520 ,
         \U1/aes_core/SB2/n2519 , \U1/aes_core/SB2/n2518 ,
         \U1/aes_core/SB2/n2517 , \U1/aes_core/SB2/n2516 ,
         \U1/aes_core/SB2/n2515 , \U1/aes_core/SB2/n2514 ,
         \U1/aes_core/SB2/n2513 , \U1/aes_core/SB2/n2512 ,
         \U1/aes_core/SB2/n2511 , \U1/aes_core/SB2/n2510 ,
         \U1/aes_core/SB2/n2509 , \U1/aes_core/SB2/n2508 ,
         \U1/aes_core/SB2/n2507 , \U1/aes_core/SB2/n2506 ,
         \U1/aes_core/SB2/n2505 , \U1/aes_core/SB2/n2504 ,
         \U1/aes_core/SB2/n2503 , \U1/aes_core/SB2/n2502 ,
         \U1/aes_core/SB2/n2501 , \U1/aes_core/SB2/n2500 ,
         \U1/aes_core/SB2/n2499 , \U1/aes_core/SB2/n2498 ,
         \U1/aes_core/SB2/n2497 , \U1/aes_core/SB2/n2496 ,
         \U1/aes_core/SB2/n2495 , \U1/aes_core/SB2/n2494 ,
         \U1/aes_core/SB2/n2493 , \U1/aes_core/SB2/n2492 ,
         \U1/aes_core/SB2/n2491 , \U1/aes_core/SB2/n2490 ,
         \U1/aes_core/SB2/n2489 , \U1/aes_core/SB2/n2488 ,
         \U1/aes_core/SB2/n2487 , \U1/aes_core/SB2/n2486 ,
         \U1/aes_core/SB2/n2485 , \U1/aes_core/SB2/n2484 ,
         \U1/aes_core/SB2/n2483 , \U1/aes_core/SB2/n2482 ,
         \U1/aes_core/SB2/n2481 , \U1/aes_core/SB2/n2480 ,
         \U1/aes_core/SB2/n2479 , \U1/aes_core/SB2/n2478 ,
         \U1/aes_core/SB2/n2477 , \U1/aes_core/SB2/n2476 ,
         \U1/aes_core/SB2/n2475 , \U1/aes_core/SB2/n2474 ,
         \U1/aes_core/SB2/n2473 , \U1/aes_core/SB2/n2472 ,
         \U1/aes_core/SB2/n2471 , \U1/aes_core/SB2/n2470 ,
         \U1/aes_core/SB2/n2469 , \U1/aes_core/SB2/n2468 ,
         \U1/aes_core/SB2/n2467 , \U1/aes_core/SB2/n2466 ,
         \U1/aes_core/SB2/n2465 , \U1/aes_core/SB2/n2464 ,
         \U1/aes_core/SB2/n2463 , \U1/aes_core/SB2/n2462 ,
         \U1/aes_core/SB2/n2461 , \U1/aes_core/SB2/n2460 ,
         \U1/aes_core/SB2/n2459 , \U1/aes_core/SB2/n2458 ,
         \U1/aes_core/SB2/n2457 , \U1/aes_core/SB2/n2456 ,
         \U1/aes_core/SB2/n2455 , \U1/aes_core/SB2/n2454 ,
         \U1/aes_core/SB2/n2453 , \U1/aes_core/SB2/n2452 ,
         \U1/aes_core/SB2/n2451 , \U1/aes_core/SB2/n2450 ,
         \U1/aes_core/SB2/n2449 , \U1/aes_core/SB2/n2448 ,
         \U1/aes_core/SB2/n2447 , \U1/aes_core/SB2/n2446 ,
         \U1/aes_core/SB2/n2445 , \U1/aes_core/SB2/n2444 ,
         \U1/aes_core/SB2/n2443 , \U1/aes_core/SB2/n2442 ,
         \U1/aes_core/SB2/n2441 , \U1/aes_core/SB2/n2440 ,
         \U1/aes_core/SB2/n2439 , \U1/aes_core/SB2/n2438 ,
         \U1/aes_core/SB2/n2437 , \U1/aes_core/SB2/n2436 ,
         \U1/aes_core/SB2/n2435 , \U1/aes_core/SB2/n2434 ,
         \U1/aes_core/SB2/n2433 , \U1/aes_core/SB2/n2432 ,
         \U1/aes_core/SB2/n2431 , \U1/aes_core/SB2/n2430 ,
         \U1/aes_core/SB2/n2429 , \U1/aes_core/SB2/n2428 ,
         \U1/aes_core/SB2/n2427 , \U1/aes_core/SB2/n2426 ,
         \U1/aes_core/SB2/n2425 , \U1/aes_core/SB2/n2424 ,
         \U1/aes_core/SB2/n2423 , \U1/aes_core/SB2/n2422 ,
         \U1/aes_core/SB2/n2421 , \U1/aes_core/SB2/n2420 ,
         \U1/aes_core/SB2/n2419 , \U1/aes_core/SB2/n2418 ,
         \U1/aes_core/SB2/n2417 , \U1/aes_core/SB2/n2416 ,
         \U1/aes_core/SB2/n2415 , \U1/aes_core/SB2/n2414 ,
         \U1/aes_core/SB2/n2413 , \U1/aes_core/SB2/n2412 ,
         \U1/aes_core/SB2/n2411 , \U1/aes_core/SB2/n2410 ,
         \U1/aes_core/SB2/n2409 , \U1/aes_core/SB2/n2408 ,
         \U1/aes_core/SB2/n2407 , \U1/aes_core/SB2/n2406 ,
         \U1/aes_core/SB2/n2405 , \U1/aes_core/SB2/n2404 ,
         \U1/aes_core/SB2/n2403 , \U1/aes_core/SB2/n2402 ,
         \U1/aes_core/SB2/n2401 , \U1/aes_core/SB2/n2400 ,
         \U1/aes_core/SB2/n2399 , \U1/aes_core/SB2/n2398 ,
         \U1/aes_core/SB2/n2397 , \U1/aes_core/SB2/n2396 ,
         \U1/aes_core/SB2/n2395 , \U1/aes_core/SB2/n2394 ,
         \U1/aes_core/SB2/n2393 , \U1/aes_core/SB2/n2392 ,
         \U1/aes_core/SB2/n2391 , \U1/aes_core/SB2/n2390 ,
         \U1/aes_core/SB2/n2389 , \U1/aes_core/SB2/n2388 ,
         \U1/aes_core/SB2/n2387 , \U1/aes_core/SB2/n2386 ,
         \U1/aes_core/SB2/n2385 , \U1/aes_core/SB2/n2384 ,
         \U1/aes_core/SB2/n2383 , \U1/aes_core/SB2/n2382 ,
         \U1/aes_core/SB2/n2381 , \U1/aes_core/SB2/n2380 ,
         \U1/aes_core/SB2/n2379 , \U1/aes_core/SB2/n2378 ,
         \U1/aes_core/SB2/n2377 , \U1/aes_core/SB2/n2376 ,
         \U1/aes_core/SB2/n2375 , \U1/aes_core/SB2/n2374 ,
         \U1/aes_core/SB2/n2373 , \U1/aes_core/SB2/n2372 ,
         \U1/aes_core/SB2/n2371 , \U1/aes_core/SB2/n2370 ,
         \U1/aes_core/SB2/n2369 , \U1/aes_core/SB2/n2368 ,
         \U1/aes_core/SB2/n2367 , \U1/aes_core/SB2/n2366 ,
         \U1/aes_core/SB2/n2365 , \U1/aes_core/SB2/n2364 ,
         \U1/aes_core/SB2/n2363 , \U1/aes_core/SB2/n2362 ,
         \U1/aes_core/SB2/n2361 , \U1/aes_core/SB2/n2360 ,
         \U1/aes_core/SB2/n2359 , \U1/aes_core/SB2/n2358 ,
         \U1/aes_core/SB2/n2357 , \U1/aes_core/SB2/n2356 ,
         \U1/aes_core/SB2/n2355 , \U1/aes_core/SB2/n2354 ,
         \U1/aes_core/SB2/n2353 , \U1/aes_core/SB2/n2352 ,
         \U1/aes_core/SB2/n2351 , \U1/aes_core/SB2/n2350 ,
         \U1/aes_core/SB2/n2349 , \U1/aes_core/SB2/n2348 ,
         \U1/aes_core/SB2/n2347 , \U1/aes_core/SB2/n2346 ,
         \U1/aes_core/SB2/n2345 , \U1/aes_core/SB2/n2344 ,
         \U1/aes_core/SB2/n2343 , \U1/aes_core/SB2/n2342 ,
         \U1/aes_core/SB2/n2341 , \U1/aes_core/SB2/n2340 ,
         \U1/aes_core/SB2/n2339 , \U1/aes_core/SB2/n2338 ,
         \U1/aes_core/SB2/n2337 , \U1/aes_core/SB2/n2336 ,
         \U1/aes_core/SB2/n2335 , \U1/aes_core/SB2/n2334 ,
         \U1/aes_core/SB2/n2333 , \U1/aes_core/SB2/n2332 ,
         \U1/aes_core/SB2/n2331 , \U1/aes_core/SB2/n2330 ,
         \U1/aes_core/SB2/n2329 , \U1/aes_core/SB2/n2328 ,
         \U1/aes_core/SB2/n2327 , \U1/aes_core/SB2/n2326 ,
         \U1/aes_core/SB2/n2325 , \U1/aes_core/SB2/n2324 ,
         \U1/aes_core/SB2/n2323 , \U1/aes_core/SB2/n2322 ,
         \U1/aes_core/SB2/n2321 , \U1/aes_core/SB2/n2320 ,
         \U1/aes_core/SB2/n2319 , \U1/aes_core/SB2/n2318 ,
         \U1/aes_core/SB2/n2317 , \U1/aes_core/SB2/n2316 ,
         \U1/aes_core/SB2/n2315 , \U1/aes_core/SB2/n2314 ,
         \U1/aes_core/SB2/n2313 , \U1/aes_core/SB2/n2312 ,
         \U1/aes_core/SB2/n2311 , \U1/aes_core/SB2/n2310 ,
         \U1/aes_core/SB2/n2309 , \U1/aes_core/SB2/n2308 ,
         \U1/aes_core/SB2/n2307 , \U1/aes_core/SB2/n2306 ,
         \U1/aes_core/SB2/n2305 , \U1/aes_core/SB2/n2304 ,
         \U1/aes_core/SB2/n2303 , \U1/aes_core/SB2/n2302 ,
         \U1/aes_core/SB2/n2301 , \U1/aes_core/SB2/n2300 ,
         \U1/aes_core/SB2/n2299 , \U1/aes_core/SB2/n2298 ,
         \U1/aes_core/SB2/n2297 , \U1/aes_core/SB2/n2296 ,
         \U1/aes_core/SB2/n2295 , \U1/aes_core/SB2/n2294 ,
         \U1/aes_core/SB2/n2293 , \U1/aes_core/SB2/n2292 ,
         \U1/aes_core/SB2/n2291 , \U1/aes_core/SB2/n2290 ,
         \U1/aes_core/SB2/n2289 , \U1/aes_core/SB2/n2288 ,
         \U1/aes_core/SB2/n2287 , \U1/aes_core/SB2/n2286 ,
         \U1/aes_core/SB2/n2285 , \U1/aes_core/SB2/n2284 ,
         \U1/aes_core/SB2/n2283 , \U1/aes_core/SB2/n2282 ,
         \U1/aes_core/SB2/n2281 , \U1/aes_core/SB2/n2280 ,
         \U1/aes_core/SB2/n2279 , \U1/aes_core/SB2/n2278 ,
         \U1/aes_core/SB2/n2277 , \U1/aes_core/SB2/n2276 ,
         \U1/aes_core/SB2/n2275 , \U1/aes_core/SB2/n2274 ,
         \U1/aes_core/SB2/n2273 , \U1/aes_core/SB2/n2272 ,
         \U1/aes_core/SB2/n2271 , \U1/aes_core/SB2/n2270 ,
         \U1/aes_core/SB2/n2269 , \U1/aes_core/SB2/n2268 ,
         \U1/aes_core/SB2/n2267 , \U1/aes_core/SB2/n2266 ,
         \U1/aes_core/SB2/n2265 , \U1/aes_core/SB2/n2264 ,
         \U1/aes_core/SB2/n2263 , \U1/aes_core/SB2/n2262 ,
         \U1/aes_core/SB2/n2261 , \U1/aes_core/SB2/n2260 ,
         \U1/aes_core/SB2/n2259 , \U1/aes_core/SB2/n2258 ,
         \U1/aes_core/SB2/n2257 , \U1/aes_core/SB2/n2256 ,
         \U1/aes_core/SB2/n2255 , \U1/aes_core/SB2/n2254 ,
         \U1/aes_core/SB2/n2253 , \U1/aes_core/SB2/n2252 ,
         \U1/aes_core/SB2/n2251 , \U1/aes_core/SB2/n2250 ,
         \U1/aes_core/SB2/n2249 , \U1/aes_core/SB2/n2248 ,
         \U1/aes_core/SB2/n2247 , \U1/aes_core/SB2/n2246 ,
         \U1/aes_core/SB2/n2245 , \U1/aes_core/SB2/n2244 ,
         \U1/aes_core/SB2/n2243 , \U1/aes_core/SB2/n2242 ,
         \U1/aes_core/SB2/n2241 , \U1/aes_core/SB2/n2240 ,
         \U1/aes_core/SB2/n2239 , \U1/aes_core/SB2/n2238 ,
         \U1/aes_core/SB2/n2237 , \U1/aes_core/SB2/n2236 ,
         \U1/aes_core/SB2/n2235 , \U1/aes_core/SB2/n2234 ,
         \U1/aes_core/SB2/n2233 , \U1/aes_core/SB2/n2232 ,
         \U1/aes_core/SB2/n2231 , \U1/aes_core/SB2/n2230 ,
         \U1/aes_core/SB2/n2229 , \U1/aes_core/SB2/n2228 ,
         \U1/aes_core/SB2/n2227 , \U1/aes_core/SB2/n2226 ,
         \U1/aes_core/SB2/n2225 , \U1/aes_core/SB2/n2224 ,
         \U1/aes_core/SB2/n2223 , \U1/aes_core/SB2/n2222 ,
         \U1/aes_core/SB2/n2221 , \U1/aes_core/SB2/n2220 ,
         \U1/aes_core/SB2/n2219 , \U1/aes_core/SB2/n2218 ,
         \U1/aes_core/SB2/n2217 , \U1/aes_core/SB2/n2216 ,
         \U1/aes_core/SB2/n2215 , \U1/aes_core/SB2/n2214 ,
         \U1/aes_core/SB2/n2213 , \U1/aes_core/SB2/n2212 ,
         \U1/aes_core/SB2/n2211 , \U1/aes_core/SB2/n2210 ,
         \U1/aes_core/SB2/n2209 , \U1/aes_core/SB2/n2208 ,
         \U1/aes_core/SB2/n2207 , \U1/aes_core/SB2/n2206 ,
         \U1/aes_core/SB2/n2205 , \U1/aes_core/SB2/n2204 ,
         \U1/aes_core/SB2/n2203 , \U1/aes_core/SB2/n2202 ,
         \U1/aes_core/SB2/n2201 , \U1/aes_core/SB2/n2200 ,
         \U1/aes_core/SB2/n2199 , \U1/aes_core/SB2/n2198 ,
         \U1/aes_core/SB2/n2197 , \U1/aes_core/SB2/n2196 ,
         \U1/aes_core/SB2/n2195 , \U1/aes_core/SB2/n2194 ,
         \U1/aes_core/SB2/n2193 , \U1/aes_core/SB2/n2192 ,
         \U1/aes_core/SB2/n2191 , \U1/aes_core/SB2/n2190 ,
         \U1/aes_core/SB2/n2189 , \U1/aes_core/SB2/n2188 ,
         \U1/aes_core/SB2/n2187 , \U1/aes_core/SB2/n2186 ,
         \U1/aes_core/SB2/n2185 , \U1/aes_core/SB2/n2184 ,
         \U1/aes_core/SB2/n2183 , \U1/aes_core/SB2/n2182 ,
         \U1/aes_core/SB2/n2181 , \U1/aes_core/SB2/n2180 ,
         \U1/aes_core/SB2/n2179 , \U1/aes_core/SB2/n2178 ,
         \U1/aes_core/SB2/n2177 , \U1/aes_core/SB2/n2176 ,
         \U1/aes_core/SB2/n2175 , \U1/aes_core/SB2/n2174 ,
         \U1/aes_core/SB2/n2173 , \U1/aes_core/SB2/n2172 ,
         \U1/aes_core/SB2/n2171 , \U1/aes_core/SB2/n2170 ,
         \U1/aes_core/SB2/n2169 , \U1/aes_core/SB2/n2168 ,
         \U1/aes_core/SB2/n2167 , \U1/aes_core/SB2/n2166 ,
         \U1/aes_core/SB2/n2165 , \U1/aes_core/SB2/n2164 ,
         \U1/aes_core/SB2/n2163 , \U1/aes_core/SB2/n2162 ,
         \U1/aes_core/SB2/n2161 , \U1/aes_core/SB2/n2160 ,
         \U1/aes_core/SB2/n2159 , \U1/aes_core/SB2/n2158 ,
         \U1/aes_core/SB2/n2157 , \U1/aes_core/SB2/n2156 ,
         \U1/aes_core/SB2/n2155 , \U1/aes_core/SB2/n2154 ,
         \U1/aes_core/SB2/n2153 , \U1/aes_core/SB2/n2152 ,
         \U1/aes_core/SB2/n2151 , \U1/aes_core/SB2/n2150 ,
         \U1/aes_core/SB2/n2149 , \U1/aes_core/SB2/n2148 ,
         \U1/aes_core/SB2/n2147 , \U1/aes_core/SB2/n2146 ,
         \U1/aes_core/SB2/n2145 , \U1/aes_core/SB2/n2144 ,
         \U1/aes_core/SB2/n2143 , \U1/aes_core/SB2/n2142 ,
         \U1/aes_core/SB2/n2141 , \U1/aes_core/SB2/n2140 ,
         \U1/aes_core/SB2/n2139 , \U1/aes_core/SB2/n2138 ,
         \U1/aes_core/SB2/n2137 , \U1/aes_core/SB2/n2136 ,
         \U1/aes_core/SB2/n2135 , \U1/aes_core/SB2/n2134 ,
         \U1/aes_core/SB2/n2133 , \U1/aes_core/SB2/n2132 ,
         \U1/aes_core/SB2/n2131 , \U1/aes_core/SB2/n2130 ,
         \U1/aes_core/SB2/n2129 , \U1/aes_core/SB2/n2128 ,
         \U1/aes_core/SB2/n2127 , \U1/aes_core/SB2/n2126 ,
         \U1/aes_core/SB2/n2125 , \U1/aes_core/SB2/n2124 ,
         \U1/aes_core/SB2/n2123 , \U1/aes_core/SB2/n2122 ,
         \U1/aes_core/SB2/n2121 , \U1/aes_core/SB2/n2120 ,
         \U1/aes_core/SB2/n2119 , \U1/aes_core/SB2/n2118 ,
         \U1/aes_core/SB2/n2117 , \U1/aes_core/SB2/n2116 ,
         \U1/aes_core/SB2/n2115 , \U1/aes_core/SB2/n2114 ,
         \U1/aes_core/SB2/n2113 , \U1/aes_core/SB2/n2112 ,
         \U1/aes_core/SB2/n2111 , \U1/aes_core/SB2/n2110 ,
         \U1/aes_core/SB2/n2109 , \U1/aes_core/SB2/n2108 ,
         \U1/aes_core/SB2/n2107 , \U1/aes_core/SB2/n2106 ,
         \U1/aes_core/SB2/n2105 , \U1/aes_core/SB2/n2104 ,
         \U1/aes_core/SB2/n2103 , \U1/aes_core/SB2/n2102 ,
         \U1/aes_core/SB2/n2101 , \U1/aes_core/SB2/n2100 ,
         \U1/aes_core/SB2/n2099 , \U1/aes_core/SB2/n2098 ,
         \U1/aes_core/SB2/n2097 , \U1/aes_core/SB2/n2096 ,
         \U1/aes_core/SB2/n2095 , \U1/aes_core/SB2/n2094 ,
         \U1/aes_core/SB2/n2093 , \U1/aes_core/SB2/n2092 ,
         \U1/aes_core/SB2/n2091 , \U1/aes_core/SB2/n2090 ,
         \U1/aes_core/SB2/n2089 , \U1/aes_core/SB2/n2088 ,
         \U1/aes_core/SB2/n2087 , \U1/aes_core/SB2/n2086 ,
         \U1/aes_core/SB2/n2085 , \U1/aes_core/SB2/n2084 ,
         \U1/aes_core/SB2/n2083 , \U1/aes_core/SB2/n2082 ,
         \U1/aes_core/SB2/n2081 , \U1/aes_core/SB2/n2080 ,
         \U1/aes_core/SB2/n2079 , \U1/aes_core/SB2/n2078 ,
         \U1/aes_core/SB2/n2077 , \U1/aes_core/SB2/n2076 ,
         \U1/aes_core/SB2/n2075 , \U1/aes_core/SB2/n2074 ,
         \U1/aes_core/SB2/n2073 , \U1/aes_core/SB2/n2072 ,
         \U1/aes_core/SB2/n2071 , \U1/aes_core/SB2/n2070 ,
         \U1/aes_core/SB2/n2069 , \U1/aes_core/SB2/n2068 ,
         \U1/aes_core/SB2/n2067 , \U1/aes_core/SB2/n2066 ,
         \U1/aes_core/SB2/n2065 , \U1/aes_core/SB2/n2064 ,
         \U1/aes_core/SB2/n2063 , \U1/aes_core/SB2/n2062 ,
         \U1/aes_core/SB2/n2061 , \U1/aes_core/SB2/n2060 ,
         \U1/aes_core/SB2/n2059 , \U1/aes_core/SB2/n2058 ,
         \U1/aes_core/SB2/n2057 , \U1/aes_core/SB2/n2056 ,
         \U1/aes_core/SB2/n2055 , \U1/aes_core/SB2/n2054 ,
         \U1/aes_core/SB2/n2053 , \U1/aes_core/SB2/n2052 ,
         \U1/aes_core/SB2/n2051 , \U1/aes_core/SB2/n2050 ,
         \U1/aes_core/SB2/n2049 , \U1/aes_core/SB2/n2048 ,
         \U1/aes_core/SB2/n2047 , \U1/aes_core/SB2/n2046 ,
         \U1/aes_core/SB2/n2045 , \U1/aes_core/SB2/n2044 ,
         \U1/aes_core/SB2/n2043 , \U1/aes_core/SB2/n2042 ,
         \U1/aes_core/SB2/n2041 , \U1/aes_core/SB2/n2040 ,
         \U1/aes_core/SB2/n2039 , \U1/aes_core/SB2/n2038 ,
         \U1/aes_core/SB2/n2037 , \U1/aes_core/SB2/n2036 ,
         \U1/aes_core/SB2/n2035 , \U1/aes_core/SB2/n2034 ,
         \U1/aes_core/SB2/n2033 , \U1/aes_core/SB2/n2032 ,
         \U1/aes_core/SB2/n2031 , \U1/aes_core/SB2/n2030 ,
         \U1/aes_core/SB2/n2029 , \U1/aes_core/SB2/n2028 ,
         \U1/aes_core/SB2/n2027 , \U1/aes_core/SB2/n2026 ,
         \U1/aes_core/SB2/n2025 , \U1/aes_core/SB2/n2024 ,
         \U1/aes_core/SB2/n2023 , \U1/aes_core/SB2/n2022 ,
         \U1/aes_core/SB2/n2021 , \U1/aes_core/SB2/n2020 ,
         \U1/aes_core/SB2/n2019 , \U1/aes_core/SB2/n2018 ,
         \U1/aes_core/SB2/n2017 , \U1/aes_core/SB2/n2016 ,
         \U1/aes_core/SB2/n2015 , \U1/aes_core/SB2/n2014 ,
         \U1/aes_core/SB2/n2013 , \U1/aes_core/SB2/n2012 ,
         \U1/aes_core/SB2/n2011 , \U1/aes_core/SB2/n2010 ,
         \U1/aes_core/SB2/n2009 , \U1/aes_core/SB2/n2008 ,
         \U1/aes_core/SB2/n2007 , \U1/aes_core/SB2/n2006 ,
         \U1/aes_core/SB2/n2005 , \U1/aes_core/SB2/n2004 ,
         \U1/aes_core/SB2/n2003 , \U1/aes_core/SB2/n2002 ,
         \U1/aes_core/SB2/n2001 , \U1/aes_core/SB2/n2000 ,
         \U1/aes_core/SB2/n1999 , \U1/aes_core/SB2/n1998 ,
         \U1/aes_core/SB2/n1997 , \U1/aes_core/SB2/n1996 ,
         \U1/aes_core/SB2/n1995 , \U1/aes_core/SB2/n1994 ,
         \U1/aes_core/SB2/n1993 , \U1/aes_core/SB2/n1992 ,
         \U1/aes_core/SB2/n1991 , \U1/aes_core/SB2/n1990 ,
         \U1/aes_core/SB2/n1989 , \U1/aes_core/SB2/n1988 ,
         \U1/aes_core/SB2/n1987 , \U1/aes_core/SB2/n1986 ,
         \U1/aes_core/SB2/n1985 , \U1/aes_core/SB2/n1984 ,
         \U1/aes_core/SB2/n1983 , \U1/aes_core/SB2/n1982 ,
         \U1/aes_core/SB2/n1981 , \U1/aes_core/SB2/n1980 ,
         \U1/aes_core/SB2/n1979 , \U1/aes_core/SB2/n1978 ,
         \U1/aes_core/SB2/n1977 , \U1/aes_core/SB2/n1976 ,
         \U1/aes_core/SB2/n1975 , \U1/aes_core/SB2/n1974 ,
         \U1/aes_core/SB2/n1973 , \U1/aes_core/SB2/n1972 ,
         \U1/aes_core/SB2/n1971 , \U1/aes_core/SB2/n1970 ,
         \U1/aes_core/SB2/n1969 , \U1/aes_core/SB2/n1968 ,
         \U1/aes_core/SB2/n1967 , \U1/aes_core/SB2/n1966 ,
         \U1/aes_core/SB2/n1965 , \U1/aes_core/SB2/n1964 ,
         \U1/aes_core/SB2/n1963 , \U1/aes_core/SB2/n1962 ,
         \U1/aes_core/SB2/n1961 , \U1/aes_core/SB2/n1960 ,
         \U1/aes_core/SB2/n1959 , \U1/aes_core/SB2/n1958 ,
         \U1/aes_core/SB2/n1957 , \U1/aes_core/SB2/n1956 ,
         \U1/aes_core/SB2/n1955 , \U1/aes_core/SB2/n1954 ,
         \U1/aes_core/SB2/n1953 , \U1/aes_core/SB2/n1952 ,
         \U1/aes_core/SB2/n1951 , \U1/aes_core/SB2/n1950 ,
         \U1/aes_core/SB2/n1949 , \U1/aes_core/SB2/n1948 ,
         \U1/aes_core/SB2/n1947 , \U1/aes_core/SB2/n1946 ,
         \U1/aes_core/SB2/n1945 , \U1/aes_core/SB2/n1944 ,
         \U1/aes_core/SB2/n1943 , \U1/aes_core/SB2/n1942 ,
         \U1/aes_core/SB2/n1941 , \U1/aes_core/SB2/n1940 ,
         \U1/aes_core/SB2/n1939 , \U1/aes_core/SB2/n1938 ,
         \U1/aes_core/SB2/n1937 , \U1/aes_core/SB2/n1936 ,
         \U1/aes_core/SB2/n1935 , \U1/aes_core/SB2/n1934 ,
         \U1/aes_core/SB2/n1933 , \U1/aes_core/SB2/n1932 ,
         \U1/aes_core/SB2/n1931 , \U1/aes_core/SB2/n1930 ,
         \U1/aes_core/SB2/n1929 , \U1/aes_core/SB2/n1928 ,
         \U1/aes_core/SB2/n1927 , \U1/aes_core/SB2/n1926 ,
         \U1/aes_core/SB2/n1925 , \U1/aes_core/SB2/n1924 ,
         \U1/aes_core/SB2/n1923 , \U1/aes_core/SB2/n1922 ,
         \U1/aes_core/SB2/n1921 , \U1/aes_core/SB2/n1920 ,
         \U1/aes_core/SB2/n1919 , \U1/aes_core/SB2/n1918 ,
         \U1/aes_core/SB2/n1917 , \U1/aes_core/SB2/n1916 ,
         \U1/aes_core/SB2/n1915 , \U1/aes_core/SB2/n1914 ,
         \U1/aes_core/SB2/n1913 , \U1/aes_core/SB2/n1912 ,
         \U1/aes_core/SB2/n1911 , \U1/aes_core/SB2/n1910 ,
         \U1/aes_core/SB2/n1909 , \U1/aes_core/SB2/n1908 ,
         \U1/aes_core/SB2/n1907 , \U1/aes_core/SB2/n1906 ,
         \U1/aes_core/SB2/n1905 , \U1/aes_core/SB2/n1904 ,
         \U1/aes_core/SB2/n1903 , \U1/aes_core/SB2/n1902 ,
         \U1/aes_core/SB2/n1901 , \U1/aes_core/SB2/n1900 ,
         \U1/aes_core/SB2/n1899 , \U1/aes_core/SB2/n1898 ,
         \U1/aes_core/SB2/n1897 , \U1/aes_core/SB2/n1896 ,
         \U1/aes_core/SB2/n1895 , \U1/aes_core/SB2/n1894 ,
         \U1/aes_core/SB2/n1893 , \U1/aes_core/SB2/n1892 ,
         \U1/aes_core/SB2/n1891 , \U1/aes_core/SB2/n1890 ,
         \U1/aes_core/SB2/n1889 , \U1/aes_core/SB2/n1888 ,
         \U1/aes_core/SB2/n1887 , \U1/aes_core/SB2/n1886 ,
         \U1/aes_core/SB2/n1885 , \U1/aes_core/SB2/n1884 ,
         \U1/aes_core/SB2/n1883 , \U1/aes_core/SB2/n1882 ,
         \U1/aes_core/SB2/n1881 , \U1/aes_core/SB2/n1880 ,
         \U1/aes_core/SB2/n1879 , \U1/aes_core/SB2/n1878 ,
         \U1/aes_core/SB2/n1877 , \U1/aes_core/SB2/n1876 ,
         \U1/aes_core/SB2/n1875 , \U1/aes_core/SB2/n1874 ,
         \U1/aes_core/SB2/n1873 , \U1/aes_core/SB2/n1872 ,
         \U1/aes_core/SB2/n1871 , \U1/aes_core/SB2/n1870 ,
         \U1/aes_core/SB2/n1869 , \U1/aes_core/SB2/n1868 ,
         \U1/aes_core/SB2/n1867 , \U1/aes_core/SB2/n1866 ,
         \U1/aes_core/SB2/n1865 , \U1/aes_core/SB2/n1864 ,
         \U1/aes_core/SB2/n1863 , \U1/aes_core/SB2/n1862 ,
         \U1/aes_core/SB2/n1861 , \U1/aes_core/SB2/n1860 ,
         \U1/aes_core/SB2/n1859 , \U1/aes_core/SB2/n1858 ,
         \U1/aes_core/SB2/n1857 , \U1/aes_core/SB2/n1856 ,
         \U1/aes_core/SB2/n1855 , \U1/aes_core/SB2/n1854 ,
         \U1/aes_core/SB2/n1853 , \U1/aes_core/SB2/n1852 ,
         \U1/aes_core/SB2/n1851 , \U1/aes_core/SB2/n1850 ,
         \U1/aes_core/SB2/n1849 , \U1/aes_core/SB2/n1848 ,
         \U1/aes_core/SB2/n1847 , \U1/aes_core/SB2/n1846 ,
         \U1/aes_core/SB2/n1845 , \U1/aes_core/SB2/n1844 ,
         \U1/aes_core/SB2/n1843 , \U1/aes_core/SB2/n1842 ,
         \U1/aes_core/SB2/n1841 , \U1/aes_core/SB2/n1840 ,
         \U1/aes_core/SB2/n1839 , \U1/aes_core/SB2/n1838 ,
         \U1/aes_core/SB2/n1837 , \U1/aes_core/SB2/n1836 ,
         \U1/aes_core/SB2/n1835 , \U1/aes_core/SB2/n1834 ,
         \U1/aes_core/SB2/n1833 , \U1/aes_core/SB2/n1832 ,
         \U1/aes_core/SB2/n1831 , \U1/aes_core/SB2/n1830 ,
         \U1/aes_core/SB2/n1829 , \U1/aes_core/SB2/n1828 ,
         \U1/aes_core/SB2/n1827 , \U1/aes_core/SB2/n1826 ,
         \U1/aes_core/SB2/n1825 , \U1/aes_core/SB2/n1824 ,
         \U1/aes_core/SB2/n1823 , \U1/aes_core/SB2/n1822 ,
         \U1/aes_core/SB2/n1821 , \U1/aes_core/SB2/n1820 ,
         \U1/aes_core/SB2/n1819 , \U1/aes_core/SB2/n1818 ,
         \U1/aes_core/SB2/n1817 , \U1/aes_core/SB2/n1816 ,
         \U1/aes_core/SB2/n1815 , \U1/aes_core/SB2/n1814 ,
         \U1/aes_core/SB2/n1813 , \U1/aes_core/SB2/n1812 ,
         \U1/aes_core/SB2/n1811 , \U1/aes_core/SB2/n1810 ,
         \U1/aes_core/SB2/n1809 , \U1/aes_core/SB2/n1808 ,
         \U1/aes_core/SB2/n1807 , \U1/aes_core/SB2/n1806 ,
         \U1/aes_core/SB2/n1805 , \U1/aes_core/SB2/n1804 ,
         \U1/aes_core/SB2/n1803 , \U1/aes_core/SB2/n1802 ,
         \U1/aes_core/SB2/n1801 , \U1/aes_core/SB2/n1800 ,
         \U1/aes_core/SB2/n1799 , \U1/aes_core/SB2/n1798 ,
         \U1/aes_core/SB2/n1797 , \U1/aes_core/SB2/n1796 ,
         \U1/aes_core/SB2/n1795 , \U1/aes_core/SB2/n1794 ,
         \U1/aes_core/SB2/n1793 , \U1/aes_core/SB2/n1792 ,
         \U1/aes_core/SB2/n1791 , \U1/aes_core/SB2/n1790 ,
         \U1/aes_core/SB2/n1789 , \U1/aes_core/SB2/n1788 ,
         \U1/aes_core/SB2/n1787 , \U1/aes_core/SB2/n1786 ,
         \U1/aes_core/SB2/n1785 , \U1/aes_core/SB2/n1784 ,
         \U1/aes_core/SB2/n1783 , \U1/aes_core/SB2/n1782 ,
         \U1/aes_core/SB2/n1781 , \U1/aes_core/SB2/n1780 ,
         \U1/aes_core/SB2/n1779 , \U1/aes_core/SB2/n1778 ,
         \U1/aes_core/SB2/n1777 , \U1/aes_core/SB2/n1776 ,
         \U1/aes_core/SB2/n1775 , \U1/aes_core/SB2/n1774 ,
         \U1/aes_core/SB2/n1773 , \U1/aes_core/SB2/n1772 ,
         \U1/aes_core/SB2/n1771 , \U1/aes_core/SB2/n1770 ,
         \U1/aes_core/SB2/n1769 , \U1/aes_core/SB2/n1768 ,
         \U1/aes_core/SB2/n1767 , \U1/aes_core/SB2/n1766 ,
         \U1/aes_core/SB2/n1765 , \U1/aes_core/SB2/n1764 ,
         \U1/aes_core/SB2/n1763 , \U1/aes_core/SB2/n1762 ,
         \U1/aes_core/SB2/n1761 , \U1/aes_core/SB2/n1760 ,
         \U1/aes_core/SB2/n1759 , \U1/aes_core/SB2/n1758 ,
         \U1/aes_core/SB2/n1757 , \U1/aes_core/SB2/n1756 ,
         \U1/aes_core/SB2/n1755 , \U1/aes_core/SB2/n1754 ,
         \U1/aes_core/SB2/n1753 , \U1/aes_core/SB2/n1752 ,
         \U1/aes_core/SB2/n1751 , \U1/aes_core/SB2/n1750 ,
         \U1/aes_core/SB2/n1749 , \U1/aes_core/SB2/n1748 ,
         \U1/aes_core/SB2/n1747 , \U1/aes_core/SB2/n1746 ,
         \U1/aes_core/SB2/n1745 , \U1/aes_core/SB2/n1744 ,
         \U1/aes_core/SB2/n1743 , \U1/aes_core/SB2/n1742 ,
         \U1/aes_core/SB2/n1741 , \U1/aes_core/SB2/n1740 ,
         \U1/aes_core/SB2/n1739 , \U1/aes_core/SB2/n1738 ,
         \U1/aes_core/SB2/n1737 , \U1/aes_core/SB2/n1736 ,
         \U1/aes_core/SB2/n1735 , \U1/aes_core/SB2/n1734 ,
         \U1/aes_core/SB2/n1733 , \U1/aes_core/SB2/n1732 ,
         \U1/aes_core/SB2/n1731 , \U1/aes_core/SB2/n1730 ,
         \U1/aes_core/SB2/n1729 , \U1/aes_core/SB2/n1728 ,
         \U1/aes_core/SB2/n1727 , \U1/aes_core/SB2/n1726 ,
         \U1/aes_core/SB2/n1725 , \U1/aes_core/SB2/n1724 ,
         \U1/aes_core/SB2/n1723 , \U1/aes_core/SB2/n1722 ,
         \U1/aes_core/SB2/n1721 , \U1/aes_core/SB2/n1720 ,
         \U1/aes_core/SB2/n1719 , \U1/aes_core/SB2/n1718 ,
         \U1/aes_core/SB2/n1717 , \U1/aes_core/SB2/n1716 ,
         \U1/aes_core/SB2/n1715 , \U1/aes_core/SB2/n1714 ,
         \U1/aes_core/SB2/n1713 , \U1/aes_core/SB2/n1712 ,
         \U1/aes_core/SB2/n1711 , \U1/aes_core/SB2/n1710 ,
         \U1/aes_core/SB2/n1709 , \U1/aes_core/SB2/n1708 ,
         \U1/aes_core/SB2/n1707 , \U1/aes_core/SB2/n1706 ,
         \U1/aes_core/SB2/n1705 , \U1/aes_core/SB2/n1704 ,
         \U1/aes_core/SB2/n1703 , \U1/aes_core/SB2/n1702 ,
         \U1/aes_core/SB2/n1701 , \U1/aes_core/SB2/n1700 ,
         \U1/aes_core/SB2/n1699 , \U1/aes_core/SB2/n1698 ,
         \U1/aes_core/SB2/n1697 , \U1/aes_core/SB2/n1696 ,
         \U1/aes_core/SB2/n1695 , \U1/aes_core/SB2/n1694 ,
         \U1/aes_core/SB2/n1693 , \U1/aes_core/SB2/n1692 ,
         \U1/aes_core/SB2/n1691 , \U1/aes_core/SB2/n1690 ,
         \U1/aes_core/SB2/n1689 , \U1/aes_core/SB2/n1688 ,
         \U1/aes_core/SB2/n1687 , \U1/aes_core/SB2/n1686 ,
         \U1/aes_core/SB2/n1685 , \U1/aes_core/SB2/n1684 ,
         \U1/aes_core/SB2/n1683 , \U1/aes_core/SB2/n1682 ,
         \U1/aes_core/SB2/n1621 , \U1/aes_core/SB2/n1218 ,
         \U1/aes_core/SB2/n1203 , \U1/aes_core/SB2/n1158 ,
         \U1/aes_core/SB2/n1030 , \U1/aes_core/SB2/n767 ,
         \U1/aes_core/SB2/n752 , \U1/aes_core/SB2/n707 ,
         \U1/aes_core/SB2/n385 , \U1/aes_core/SB3/n3353 ,
         \U1/aes_core/SB3/n3352 , \U1/aes_core/SB3/n3351 ,
         \U1/aes_core/SB3/n3350 , \U1/aes_core/SB3/n3349 ,
         \U1/aes_core/SB3/n3348 , \U1/aes_core/SB3/n3347 ,
         \U1/aes_core/SB3/n3346 , \U1/aes_core/SB3/n3345 ,
         \U1/aes_core/SB3/n3344 , \U1/aes_core/SB3/n3343 ,
         \U1/aes_core/SB3/n3342 , \U1/aes_core/SB3/n3341 ,
         \U1/aes_core/SB3/n3340 , \U1/aes_core/SB3/n3339 ,
         \U1/aes_core/SB3/n3338 , \U1/aes_core/SB3/n3337 ,
         \U1/aes_core/SB3/n3336 , \U1/aes_core/SB3/n3335 ,
         \U1/aes_core/SB3/n3334 , \U1/aes_core/SB3/n3333 ,
         \U1/aes_core/SB3/n3332 , \U1/aes_core/SB3/n3331 ,
         \U1/aes_core/SB3/n3330 , \U1/aes_core/SB3/n3329 ,
         \U1/aes_core/SB3/n3328 , \U1/aes_core/SB3/n3327 ,
         \U1/aes_core/SB3/n3326 , \U1/aes_core/SB3/n3325 ,
         \U1/aes_core/SB3/n3324 , \U1/aes_core/SB3/n3323 ,
         \U1/aes_core/SB3/n3322 , \U1/aes_core/SB3/n3321 ,
         \U1/aes_core/SB3/n3320 , \U1/aes_core/SB3/n3319 ,
         \U1/aes_core/SB3/n3318 , \U1/aes_core/SB3/n3317 ,
         \U1/aes_core/SB3/n3316 , \U1/aes_core/SB3/n3315 ,
         \U1/aes_core/SB3/n3314 , \U1/aes_core/SB3/n3313 ,
         \U1/aes_core/SB3/n3312 , \U1/aes_core/SB3/n3311 ,
         \U1/aes_core/SB3/n3310 , \U1/aes_core/SB3/n3309 ,
         \U1/aes_core/SB3/n3308 , \U1/aes_core/SB3/n3307 ,
         \U1/aes_core/SB3/n3306 , \U1/aes_core/SB3/n3305 ,
         \U1/aes_core/SB3/n3304 , \U1/aes_core/SB3/n3303 ,
         \U1/aes_core/SB3/n3302 , \U1/aes_core/SB3/n3301 ,
         \U1/aes_core/SB3/n3300 , \U1/aes_core/SB3/n3299 ,
         \U1/aes_core/SB3/n3298 , \U1/aes_core/SB3/n3297 ,
         \U1/aes_core/SB3/n3296 , \U1/aes_core/SB3/n3295 ,
         \U1/aes_core/SB3/n3294 , \U1/aes_core/SB3/n3293 ,
         \U1/aes_core/SB3/n3292 , \U1/aes_core/SB3/n3291 ,
         \U1/aes_core/SB3/n3290 , \U1/aes_core/SB3/n3289 ,
         \U1/aes_core/SB3/n3288 , \U1/aes_core/SB3/n3287 ,
         \U1/aes_core/SB3/n3286 , \U1/aes_core/SB3/n3285 ,
         \U1/aes_core/SB3/n3284 , \U1/aes_core/SB3/n3283 ,
         \U1/aes_core/SB3/n3282 , \U1/aes_core/SB3/n3281 ,
         \U1/aes_core/SB3/n3280 , \U1/aes_core/SB3/n3279 ,
         \U1/aes_core/SB3/n3278 , \U1/aes_core/SB3/n3277 ,
         \U1/aes_core/SB3/n3276 , \U1/aes_core/SB3/n3275 ,
         \U1/aes_core/SB3/n3274 , \U1/aes_core/SB3/n3273 ,
         \U1/aes_core/SB3/n3272 , \U1/aes_core/SB3/n3271 ,
         \U1/aes_core/SB3/n3270 , \U1/aes_core/SB3/n3269 ,
         \U1/aes_core/SB3/n3268 , \U1/aes_core/SB3/n3267 ,
         \U1/aes_core/SB3/n3266 , \U1/aes_core/SB3/n3265 ,
         \U1/aes_core/SB3/n3264 , \U1/aes_core/SB3/n3263 ,
         \U1/aes_core/SB3/n3262 , \U1/aes_core/SB3/n3261 ,
         \U1/aes_core/SB3/n3260 , \U1/aes_core/SB3/n3259 ,
         \U1/aes_core/SB3/n3258 , \U1/aes_core/SB3/n3257 ,
         \U1/aes_core/SB3/n3256 , \U1/aes_core/SB3/n3255 ,
         \U1/aes_core/SB3/n3254 , \U1/aes_core/SB3/n3253 ,
         \U1/aes_core/SB3/n3252 , \U1/aes_core/SB3/n3251 ,
         \U1/aes_core/SB3/n3250 , \U1/aes_core/SB3/n3249 ,
         \U1/aes_core/SB3/n3248 , \U1/aes_core/SB3/n3247 ,
         \U1/aes_core/SB3/n3246 , \U1/aes_core/SB3/n3245 ,
         \U1/aes_core/SB3/n3244 , \U1/aes_core/SB3/n3243 ,
         \U1/aes_core/SB3/n3242 , \U1/aes_core/SB3/n3241 ,
         \U1/aes_core/SB3/n3240 , \U1/aes_core/SB3/n3239 ,
         \U1/aes_core/SB3/n3238 , \U1/aes_core/SB3/n3237 ,
         \U1/aes_core/SB3/n3236 , \U1/aes_core/SB3/n3235 ,
         \U1/aes_core/SB3/n3234 , \U1/aes_core/SB3/n3233 ,
         \U1/aes_core/SB3/n3232 , \U1/aes_core/SB3/n3231 ,
         \U1/aes_core/SB3/n3230 , \U1/aes_core/SB3/n3229 ,
         \U1/aes_core/SB3/n3228 , \U1/aes_core/SB3/n3227 ,
         \U1/aes_core/SB3/n3226 , \U1/aes_core/SB3/n3225 ,
         \U1/aes_core/SB3/n3224 , \U1/aes_core/SB3/n3223 ,
         \U1/aes_core/SB3/n3222 , \U1/aes_core/SB3/n3221 ,
         \U1/aes_core/SB3/n3220 , \U1/aes_core/SB3/n3219 ,
         \U1/aes_core/SB3/n3218 , \U1/aes_core/SB3/n3217 ,
         \U1/aes_core/SB3/n3216 , \U1/aes_core/SB3/n3215 ,
         \U1/aes_core/SB3/n3214 , \U1/aes_core/SB3/n3213 ,
         \U1/aes_core/SB3/n3212 , \U1/aes_core/SB3/n3211 ,
         \U1/aes_core/SB3/n3210 , \U1/aes_core/SB3/n3209 ,
         \U1/aes_core/SB3/n3208 , \U1/aes_core/SB3/n3207 ,
         \U1/aes_core/SB3/n3206 , \U1/aes_core/SB3/n3205 ,
         \U1/aes_core/SB3/n3204 , \U1/aes_core/SB3/n3203 ,
         \U1/aes_core/SB3/n3202 , \U1/aes_core/SB3/n3201 ,
         \U1/aes_core/SB3/n3200 , \U1/aes_core/SB3/n3199 ,
         \U1/aes_core/SB3/n3198 , \U1/aes_core/SB3/n3197 ,
         \U1/aes_core/SB3/n3196 , \U1/aes_core/SB3/n3195 ,
         \U1/aes_core/SB3/n3194 , \U1/aes_core/SB3/n3193 ,
         \U1/aes_core/SB3/n3192 , \U1/aes_core/SB3/n3191 ,
         \U1/aes_core/SB3/n3190 , \U1/aes_core/SB3/n3189 ,
         \U1/aes_core/SB3/n3188 , \U1/aes_core/SB3/n3187 ,
         \U1/aes_core/SB3/n3186 , \U1/aes_core/SB3/n3185 ,
         \U1/aes_core/SB3/n3184 , \U1/aes_core/SB3/n3183 ,
         \U1/aes_core/SB3/n3182 , \U1/aes_core/SB3/n3181 ,
         \U1/aes_core/SB3/n3180 , \U1/aes_core/SB3/n3179 ,
         \U1/aes_core/SB3/n3178 , \U1/aes_core/SB3/n3177 ,
         \U1/aes_core/SB3/n3176 , \U1/aes_core/SB3/n3175 ,
         \U1/aes_core/SB3/n3174 , \U1/aes_core/SB3/n3173 ,
         \U1/aes_core/SB3/n3172 , \U1/aes_core/SB3/n3171 ,
         \U1/aes_core/SB3/n3170 , \U1/aes_core/SB3/n3169 ,
         \U1/aes_core/SB3/n3168 , \U1/aes_core/SB3/n3167 ,
         \U1/aes_core/SB3/n3166 , \U1/aes_core/SB3/n3165 ,
         \U1/aes_core/SB3/n3164 , \U1/aes_core/SB3/n3163 ,
         \U1/aes_core/SB3/n3162 , \U1/aes_core/SB3/n3161 ,
         \U1/aes_core/SB3/n3160 , \U1/aes_core/SB3/n3159 ,
         \U1/aes_core/SB3/n3158 , \U1/aes_core/SB3/n3157 ,
         \U1/aes_core/SB3/n3156 , \U1/aes_core/SB3/n3155 ,
         \U1/aes_core/SB3/n3154 , \U1/aes_core/SB3/n3153 ,
         \U1/aes_core/SB3/n3152 , \U1/aes_core/SB3/n3151 ,
         \U1/aes_core/SB3/n3150 , \U1/aes_core/SB3/n3149 ,
         \U1/aes_core/SB3/n3148 , \U1/aes_core/SB3/n3147 ,
         \U1/aes_core/SB3/n3146 , \U1/aes_core/SB3/n3145 ,
         \U1/aes_core/SB3/n3144 , \U1/aes_core/SB3/n3143 ,
         \U1/aes_core/SB3/n3142 , \U1/aes_core/SB3/n3141 ,
         \U1/aes_core/SB3/n3140 , \U1/aes_core/SB3/n3139 ,
         \U1/aes_core/SB3/n3138 , \U1/aes_core/SB3/n3137 ,
         \U1/aes_core/SB3/n3136 , \U1/aes_core/SB3/n3135 ,
         \U1/aes_core/SB3/n3134 , \U1/aes_core/SB3/n3133 ,
         \U1/aes_core/SB3/n3132 , \U1/aes_core/SB3/n3131 ,
         \U1/aes_core/SB3/n3130 , \U1/aes_core/SB3/n3129 ,
         \U1/aes_core/SB3/n3128 , \U1/aes_core/SB3/n3127 ,
         \U1/aes_core/SB3/n3126 , \U1/aes_core/SB3/n3125 ,
         \U1/aes_core/SB3/n3124 , \U1/aes_core/SB3/n3123 ,
         \U1/aes_core/SB3/n3122 , \U1/aes_core/SB3/n3121 ,
         \U1/aes_core/SB3/n3120 , \U1/aes_core/SB3/n3119 ,
         \U1/aes_core/SB3/n3118 , \U1/aes_core/SB3/n3117 ,
         \U1/aes_core/SB3/n3116 , \U1/aes_core/SB3/n3115 ,
         \U1/aes_core/SB3/n3114 , \U1/aes_core/SB3/n3113 ,
         \U1/aes_core/SB3/n3112 , \U1/aes_core/SB3/n3111 ,
         \U1/aes_core/SB3/n3110 , \U1/aes_core/SB3/n3109 ,
         \U1/aes_core/SB3/n3108 , \U1/aes_core/SB3/n3107 ,
         \U1/aes_core/SB3/n3106 , \U1/aes_core/SB3/n3105 ,
         \U1/aes_core/SB3/n3104 , \U1/aes_core/SB3/n3103 ,
         \U1/aes_core/SB3/n3102 , \U1/aes_core/SB3/n3101 ,
         \U1/aes_core/SB3/n3100 , \U1/aes_core/SB3/n3099 ,
         \U1/aes_core/SB3/n3098 , \U1/aes_core/SB3/n3097 ,
         \U1/aes_core/SB3/n3096 , \U1/aes_core/SB3/n3095 ,
         \U1/aes_core/SB3/n3094 , \U1/aes_core/SB3/n3093 ,
         \U1/aes_core/SB3/n3092 , \U1/aes_core/SB3/n3091 ,
         \U1/aes_core/SB3/n3090 , \U1/aes_core/SB3/n3089 ,
         \U1/aes_core/SB3/n3088 , \U1/aes_core/SB3/n3087 ,
         \U1/aes_core/SB3/n3086 , \U1/aes_core/SB3/n3085 ,
         \U1/aes_core/SB3/n3084 , \U1/aes_core/SB3/n3083 ,
         \U1/aes_core/SB3/n3082 , \U1/aes_core/SB3/n3081 ,
         \U1/aes_core/SB3/n3080 , \U1/aes_core/SB3/n3079 ,
         \U1/aes_core/SB3/n3078 , \U1/aes_core/SB3/n3077 ,
         \U1/aes_core/SB3/n3076 , \U1/aes_core/SB3/n3075 ,
         \U1/aes_core/SB3/n3074 , \U1/aes_core/SB3/n3073 ,
         \U1/aes_core/SB3/n3072 , \U1/aes_core/SB3/n3071 ,
         \U1/aes_core/SB3/n3070 , \U1/aes_core/SB3/n3069 ,
         \U1/aes_core/SB3/n3068 , \U1/aes_core/SB3/n3067 ,
         \U1/aes_core/SB3/n3066 , \U1/aes_core/SB3/n3065 ,
         \U1/aes_core/SB3/n3064 , \U1/aes_core/SB3/n3063 ,
         \U1/aes_core/SB3/n3062 , \U1/aes_core/SB3/n3061 ,
         \U1/aes_core/SB3/n3060 , \U1/aes_core/SB3/n3059 ,
         \U1/aes_core/SB3/n3058 , \U1/aes_core/SB3/n3057 ,
         \U1/aes_core/SB3/n3056 , \U1/aes_core/SB3/n3055 ,
         \U1/aes_core/SB3/n3054 , \U1/aes_core/SB3/n3053 ,
         \U1/aes_core/SB3/n3052 , \U1/aes_core/SB3/n3051 ,
         \U1/aes_core/SB3/n3050 , \U1/aes_core/SB3/n3049 ,
         \U1/aes_core/SB3/n3048 , \U1/aes_core/SB3/n3047 ,
         \U1/aes_core/SB3/n3046 , \U1/aes_core/SB3/n3045 ,
         \U1/aes_core/SB3/n3044 , \U1/aes_core/SB3/n3043 ,
         \U1/aes_core/SB3/n3042 , \U1/aes_core/SB3/n3041 ,
         \U1/aes_core/SB3/n3040 , \U1/aes_core/SB3/n3039 ,
         \U1/aes_core/SB3/n3038 , \U1/aes_core/SB3/n3037 ,
         \U1/aes_core/SB3/n3036 , \U1/aes_core/SB3/n3035 ,
         \U1/aes_core/SB3/n3034 , \U1/aes_core/SB3/n3033 ,
         \U1/aes_core/SB3/n3032 , \U1/aes_core/SB3/n3031 ,
         \U1/aes_core/SB3/n3030 , \U1/aes_core/SB3/n3029 ,
         \U1/aes_core/SB3/n3028 , \U1/aes_core/SB3/n3027 ,
         \U1/aes_core/SB3/n3026 , \U1/aes_core/SB3/n3025 ,
         \U1/aes_core/SB3/n3024 , \U1/aes_core/SB3/n3023 ,
         \U1/aes_core/SB3/n3022 , \U1/aes_core/SB3/n3021 ,
         \U1/aes_core/SB3/n3020 , \U1/aes_core/SB3/n3019 ,
         \U1/aes_core/SB3/n3018 , \U1/aes_core/SB3/n3017 ,
         \U1/aes_core/SB3/n3016 , \U1/aes_core/SB3/n3015 ,
         \U1/aes_core/SB3/n3014 , \U1/aes_core/SB3/n3013 ,
         \U1/aes_core/SB3/n3012 , \U1/aes_core/SB3/n3011 ,
         \U1/aes_core/SB3/n3010 , \U1/aes_core/SB3/n3009 ,
         \U1/aes_core/SB3/n3008 , \U1/aes_core/SB3/n3007 ,
         \U1/aes_core/SB3/n3006 , \U1/aes_core/SB3/n3005 ,
         \U1/aes_core/SB3/n3004 , \U1/aes_core/SB3/n3003 ,
         \U1/aes_core/SB3/n3002 , \U1/aes_core/SB3/n3001 ,
         \U1/aes_core/SB3/n3000 , \U1/aes_core/SB3/n2999 ,
         \U1/aes_core/SB3/n2998 , \U1/aes_core/SB3/n2997 ,
         \U1/aes_core/SB3/n2996 , \U1/aes_core/SB3/n2995 ,
         \U1/aes_core/SB3/n2994 , \U1/aes_core/SB3/n2993 ,
         \U1/aes_core/SB3/n2992 , \U1/aes_core/SB3/n2991 ,
         \U1/aes_core/SB3/n2990 , \U1/aes_core/SB3/n2989 ,
         \U1/aes_core/SB3/n2988 , \U1/aes_core/SB3/n2987 ,
         \U1/aes_core/SB3/n2986 , \U1/aes_core/SB3/n2985 ,
         \U1/aes_core/SB3/n2984 , \U1/aes_core/SB3/n2983 ,
         \U1/aes_core/SB3/n2982 , \U1/aes_core/SB3/n2981 ,
         \U1/aes_core/SB3/n2980 , \U1/aes_core/SB3/n2979 ,
         \U1/aes_core/SB3/n2978 , \U1/aes_core/SB3/n2977 ,
         \U1/aes_core/SB3/n2976 , \U1/aes_core/SB3/n2975 ,
         \U1/aes_core/SB3/n2974 , \U1/aes_core/SB3/n2973 ,
         \U1/aes_core/SB3/n2972 , \U1/aes_core/SB3/n2971 ,
         \U1/aes_core/SB3/n2970 , \U1/aes_core/SB3/n2969 ,
         \U1/aes_core/SB3/n2968 , \U1/aes_core/SB3/n2967 ,
         \U1/aes_core/SB3/n2966 , \U1/aes_core/SB3/n2965 ,
         \U1/aes_core/SB3/n2964 , \U1/aes_core/SB3/n2963 ,
         \U1/aes_core/SB3/n2962 , \U1/aes_core/SB3/n2961 ,
         \U1/aes_core/SB3/n2960 , \U1/aes_core/SB3/n2959 ,
         \U1/aes_core/SB3/n2958 , \U1/aes_core/SB3/n2957 ,
         \U1/aes_core/SB3/n2956 , \U1/aes_core/SB3/n2955 ,
         \U1/aes_core/SB3/n2954 , \U1/aes_core/SB3/n2953 ,
         \U1/aes_core/SB3/n2952 , \U1/aes_core/SB3/n2951 ,
         \U1/aes_core/SB3/n2950 , \U1/aes_core/SB3/n2949 ,
         \U1/aes_core/SB3/n2948 , \U1/aes_core/SB3/n2947 ,
         \U1/aes_core/SB3/n2946 , \U1/aes_core/SB3/n2945 ,
         \U1/aes_core/SB3/n2944 , \U1/aes_core/SB3/n2943 ,
         \U1/aes_core/SB3/n2942 , \U1/aes_core/SB3/n2941 ,
         \U1/aes_core/SB3/n2940 , \U1/aes_core/SB3/n2939 ,
         \U1/aes_core/SB3/n2938 , \U1/aes_core/SB3/n2937 ,
         \U1/aes_core/SB3/n2936 , \U1/aes_core/SB3/n2935 ,
         \U1/aes_core/SB3/n2934 , \U1/aes_core/SB3/n2933 ,
         \U1/aes_core/SB3/n2932 , \U1/aes_core/SB3/n2931 ,
         \U1/aes_core/SB3/n2930 , \U1/aes_core/SB3/n2929 ,
         \U1/aes_core/SB3/n2928 , \U1/aes_core/SB3/n2927 ,
         \U1/aes_core/SB3/n2926 , \U1/aes_core/SB3/n2925 ,
         \U1/aes_core/SB3/n2924 , \U1/aes_core/SB3/n2923 ,
         \U1/aes_core/SB3/n2922 , \U1/aes_core/SB3/n2921 ,
         \U1/aes_core/SB3/n2920 , \U1/aes_core/SB3/n2919 ,
         \U1/aes_core/SB3/n2918 , \U1/aes_core/SB3/n2917 ,
         \U1/aes_core/SB3/n2916 , \U1/aes_core/SB3/n2915 ,
         \U1/aes_core/SB3/n2914 , \U1/aes_core/SB3/n2913 ,
         \U1/aes_core/SB3/n2912 , \U1/aes_core/SB3/n2911 ,
         \U1/aes_core/SB3/n2910 , \U1/aes_core/SB3/n2909 ,
         \U1/aes_core/SB3/n2908 , \U1/aes_core/SB3/n2907 ,
         \U1/aes_core/SB3/n2906 , \U1/aes_core/SB3/n2905 ,
         \U1/aes_core/SB3/n2904 , \U1/aes_core/SB3/n2903 ,
         \U1/aes_core/SB3/n2902 , \U1/aes_core/SB3/n2901 ,
         \U1/aes_core/SB3/n2900 , \U1/aes_core/SB3/n2899 ,
         \U1/aes_core/SB3/n2898 , \U1/aes_core/SB3/n2897 ,
         \U1/aes_core/SB3/n2896 , \U1/aes_core/SB3/n2895 ,
         \U1/aes_core/SB3/n2894 , \U1/aes_core/SB3/n2893 ,
         \U1/aes_core/SB3/n2892 , \U1/aes_core/SB3/n2891 ,
         \U1/aes_core/SB3/n2890 , \U1/aes_core/SB3/n2889 ,
         \U1/aes_core/SB3/n2888 , \U1/aes_core/SB3/n2887 ,
         \U1/aes_core/SB3/n2886 , \U1/aes_core/SB3/n2885 ,
         \U1/aes_core/SB3/n2884 , \U1/aes_core/SB3/n2883 ,
         \U1/aes_core/SB3/n2882 , \U1/aes_core/SB3/n2881 ,
         \U1/aes_core/SB3/n2880 , \U1/aes_core/SB3/n2879 ,
         \U1/aes_core/SB3/n2878 , \U1/aes_core/SB3/n2877 ,
         \U1/aes_core/SB3/n2876 , \U1/aes_core/SB3/n2875 ,
         \U1/aes_core/SB3/n2874 , \U1/aes_core/SB3/n2873 ,
         \U1/aes_core/SB3/n2872 , \U1/aes_core/SB3/n2871 ,
         \U1/aes_core/SB3/n2870 , \U1/aes_core/SB3/n2869 ,
         \U1/aes_core/SB3/n2868 , \U1/aes_core/SB3/n2867 ,
         \U1/aes_core/SB3/n2866 , \U1/aes_core/SB3/n2865 ,
         \U1/aes_core/SB3/n2864 , \U1/aes_core/SB3/n2863 ,
         \U1/aes_core/SB3/n2862 , \U1/aes_core/SB3/n2861 ,
         \U1/aes_core/SB3/n2860 , \U1/aes_core/SB3/n2859 ,
         \U1/aes_core/SB3/n2858 , \U1/aes_core/SB3/n2857 ,
         \U1/aes_core/SB3/n2856 , \U1/aes_core/SB3/n2855 ,
         \U1/aes_core/SB3/n2854 , \U1/aes_core/SB3/n2853 ,
         \U1/aes_core/SB3/n2852 , \U1/aes_core/SB3/n2851 ,
         \U1/aes_core/SB3/n2850 , \U1/aes_core/SB3/n2849 ,
         \U1/aes_core/SB3/n2848 , \U1/aes_core/SB3/n2847 ,
         \U1/aes_core/SB3/n2846 , \U1/aes_core/SB3/n2845 ,
         \U1/aes_core/SB3/n2844 , \U1/aes_core/SB3/n2843 ,
         \U1/aes_core/SB3/n2842 , \U1/aes_core/SB3/n2841 ,
         \U1/aes_core/SB3/n2840 , \U1/aes_core/SB3/n2839 ,
         \U1/aes_core/SB3/n2838 , \U1/aes_core/SB3/n2837 ,
         \U1/aes_core/SB3/n2836 , \U1/aes_core/SB3/n2835 ,
         \U1/aes_core/SB3/n2834 , \U1/aes_core/SB3/n2833 ,
         \U1/aes_core/SB3/n2832 , \U1/aes_core/SB3/n2831 ,
         \U1/aes_core/SB3/n2830 , \U1/aes_core/SB3/n2829 ,
         \U1/aes_core/SB3/n2828 , \U1/aes_core/SB3/n2827 ,
         \U1/aes_core/SB3/n2826 , \U1/aes_core/SB3/n2825 ,
         \U1/aes_core/SB3/n2824 , \U1/aes_core/SB3/n2823 ,
         \U1/aes_core/SB3/n2822 , \U1/aes_core/SB3/n2821 ,
         \U1/aes_core/SB3/n2820 , \U1/aes_core/SB3/n2819 ,
         \U1/aes_core/SB3/n2818 , \U1/aes_core/SB3/n2817 ,
         \U1/aes_core/SB3/n2816 , \U1/aes_core/SB3/n2815 ,
         \U1/aes_core/SB3/n2814 , \U1/aes_core/SB3/n2813 ,
         \U1/aes_core/SB3/n2812 , \U1/aes_core/SB3/n2811 ,
         \U1/aes_core/SB3/n2810 , \U1/aes_core/SB3/n2809 ,
         \U1/aes_core/SB3/n2808 , \U1/aes_core/SB3/n2807 ,
         \U1/aes_core/SB3/n2806 , \U1/aes_core/SB3/n2805 ,
         \U1/aes_core/SB3/n2804 , \U1/aes_core/SB3/n2803 ,
         \U1/aes_core/SB3/n2802 , \U1/aes_core/SB3/n2801 ,
         \U1/aes_core/SB3/n2800 , \U1/aes_core/SB3/n2799 ,
         \U1/aes_core/SB3/n2798 , \U1/aes_core/SB3/n2797 ,
         \U1/aes_core/SB3/n2796 , \U1/aes_core/SB3/n2795 ,
         \U1/aes_core/SB3/n2794 , \U1/aes_core/SB3/n2793 ,
         \U1/aes_core/SB3/n2792 , \U1/aes_core/SB3/n2791 ,
         \U1/aes_core/SB3/n2790 , \U1/aes_core/SB3/n2789 ,
         \U1/aes_core/SB3/n2788 , \U1/aes_core/SB3/n2787 ,
         \U1/aes_core/SB3/n2786 , \U1/aes_core/SB3/n2785 ,
         \U1/aes_core/SB3/n2784 , \U1/aes_core/SB3/n2783 ,
         \U1/aes_core/SB3/n2782 , \U1/aes_core/SB3/n2781 ,
         \U1/aes_core/SB3/n2780 , \U1/aes_core/SB3/n2779 ,
         \U1/aes_core/SB3/n2778 , \U1/aes_core/SB3/n2777 ,
         \U1/aes_core/SB3/n2776 , \U1/aes_core/SB3/n2775 ,
         \U1/aes_core/SB3/n2774 , \U1/aes_core/SB3/n2773 ,
         \U1/aes_core/SB3/n2772 , \U1/aes_core/SB3/n2771 ,
         \U1/aes_core/SB3/n2770 , \U1/aes_core/SB3/n2769 ,
         \U1/aes_core/SB3/n2768 , \U1/aes_core/SB3/n2767 ,
         \U1/aes_core/SB3/n2766 , \U1/aes_core/SB3/n2765 ,
         \U1/aes_core/SB3/n2764 , \U1/aes_core/SB3/n2763 ,
         \U1/aes_core/SB3/n2762 , \U1/aes_core/SB3/n2761 ,
         \U1/aes_core/SB3/n2760 , \U1/aes_core/SB3/n2759 ,
         \U1/aes_core/SB3/n2758 , \U1/aes_core/SB3/n2757 ,
         \U1/aes_core/SB3/n2756 , \U1/aes_core/SB3/n2755 ,
         \U1/aes_core/SB3/n2754 , \U1/aes_core/SB3/n2753 ,
         \U1/aes_core/SB3/n2752 , \U1/aes_core/SB3/n2751 ,
         \U1/aes_core/SB3/n2750 , \U1/aes_core/SB3/n2749 ,
         \U1/aes_core/SB3/n2748 , \U1/aes_core/SB3/n2747 ,
         \U1/aes_core/SB3/n2746 , \U1/aes_core/SB3/n2745 ,
         \U1/aes_core/SB3/n2744 , \U1/aes_core/SB3/n2743 ,
         \U1/aes_core/SB3/n2742 , \U1/aes_core/SB3/n2741 ,
         \U1/aes_core/SB3/n2740 , \U1/aes_core/SB3/n2739 ,
         \U1/aes_core/SB3/n2738 , \U1/aes_core/SB3/n2737 ,
         \U1/aes_core/SB3/n2736 , \U1/aes_core/SB3/n2735 ,
         \U1/aes_core/SB3/n2734 , \U1/aes_core/SB3/n2733 ,
         \U1/aes_core/SB3/n2732 , \U1/aes_core/SB3/n2731 ,
         \U1/aes_core/SB3/n2730 , \U1/aes_core/SB3/n2729 ,
         \U1/aes_core/SB3/n2728 , \U1/aes_core/SB3/n2727 ,
         \U1/aes_core/SB3/n2726 , \U1/aes_core/SB3/n2725 ,
         \U1/aes_core/SB3/n2724 , \U1/aes_core/SB3/n2723 ,
         \U1/aes_core/SB3/n2722 , \U1/aes_core/SB3/n2721 ,
         \U1/aes_core/SB3/n2720 , \U1/aes_core/SB3/n2719 ,
         \U1/aes_core/SB3/n2718 , \U1/aes_core/SB3/n2717 ,
         \U1/aes_core/SB3/n2716 , \U1/aes_core/SB3/n2715 ,
         \U1/aes_core/SB3/n2714 , \U1/aes_core/SB3/n2713 ,
         \U1/aes_core/SB3/n2712 , \U1/aes_core/SB3/n2711 ,
         \U1/aes_core/SB3/n2710 , \U1/aes_core/SB3/n2709 ,
         \U1/aes_core/SB3/n2708 , \U1/aes_core/SB3/n2707 ,
         \U1/aes_core/SB3/n2706 , \U1/aes_core/SB3/n2705 ,
         \U1/aes_core/SB3/n2704 , \U1/aes_core/SB3/n2703 ,
         \U1/aes_core/SB3/n2702 , \U1/aes_core/SB3/n2701 ,
         \U1/aes_core/SB3/n2700 , \U1/aes_core/SB3/n2699 ,
         \U1/aes_core/SB3/n2698 , \U1/aes_core/SB3/n2697 ,
         \U1/aes_core/SB3/n2696 , \U1/aes_core/SB3/n2695 ,
         \U1/aes_core/SB3/n2694 , \U1/aes_core/SB3/n2693 ,
         \U1/aes_core/SB3/n2692 , \U1/aes_core/SB3/n2691 ,
         \U1/aes_core/SB3/n2690 , \U1/aes_core/SB3/n2689 ,
         \U1/aes_core/SB3/n2688 , \U1/aes_core/SB3/n2687 ,
         \U1/aes_core/SB3/n2686 , \U1/aes_core/SB3/n2685 ,
         \U1/aes_core/SB3/n2684 , \U1/aes_core/SB3/n2683 ,
         \U1/aes_core/SB3/n2682 , \U1/aes_core/SB3/n2681 ,
         \U1/aes_core/SB3/n2680 , \U1/aes_core/SB3/n2679 ,
         \U1/aes_core/SB3/n2678 , \U1/aes_core/SB3/n2677 ,
         \U1/aes_core/SB3/n2676 , \U1/aes_core/SB3/n2675 ,
         \U1/aes_core/SB3/n2674 , \U1/aes_core/SB3/n2673 ,
         \U1/aes_core/SB3/n2672 , \U1/aes_core/SB3/n2671 ,
         \U1/aes_core/SB3/n2670 , \U1/aes_core/SB3/n2669 ,
         \U1/aes_core/SB3/n2668 , \U1/aes_core/SB3/n2667 ,
         \U1/aes_core/SB3/n2666 , \U1/aes_core/SB3/n2665 ,
         \U1/aes_core/SB3/n2664 , \U1/aes_core/SB3/n2663 ,
         \U1/aes_core/SB3/n2662 , \U1/aes_core/SB3/n2661 ,
         \U1/aes_core/SB3/n2660 , \U1/aes_core/SB3/n2659 ,
         \U1/aes_core/SB3/n2658 , \U1/aes_core/SB3/n2657 ,
         \U1/aes_core/SB3/n2656 , \U1/aes_core/SB3/n2655 ,
         \U1/aes_core/SB3/n2654 , \U1/aes_core/SB3/n2653 ,
         \U1/aes_core/SB3/n2652 , \U1/aes_core/SB3/n2651 ,
         \U1/aes_core/SB3/n2650 , \U1/aes_core/SB3/n2649 ,
         \U1/aes_core/SB3/n2648 , \U1/aes_core/SB3/n2647 ,
         \U1/aes_core/SB3/n2646 , \U1/aes_core/SB3/n2645 ,
         \U1/aes_core/SB3/n2644 , \U1/aes_core/SB3/n2643 ,
         \U1/aes_core/SB3/n2642 , \U1/aes_core/SB3/n2641 ,
         \U1/aes_core/SB3/n2640 , \U1/aes_core/SB3/n2639 ,
         \U1/aes_core/SB3/n2638 , \U1/aes_core/SB3/n2637 ,
         \U1/aes_core/SB3/n2636 , \U1/aes_core/SB3/n2635 ,
         \U1/aes_core/SB3/n2634 , \U1/aes_core/SB3/n2633 ,
         \U1/aes_core/SB3/n2632 , \U1/aes_core/SB3/n2631 ,
         \U1/aes_core/SB3/n2630 , \U1/aes_core/SB3/n2629 ,
         \U1/aes_core/SB3/n2628 , \U1/aes_core/SB3/n2627 ,
         \U1/aes_core/SB3/n2626 , \U1/aes_core/SB3/n2625 ,
         \U1/aes_core/SB3/n2624 , \U1/aes_core/SB3/n2623 ,
         \U1/aes_core/SB3/n2622 , \U1/aes_core/SB3/n2621 ,
         \U1/aes_core/SB3/n2620 , \U1/aes_core/SB3/n2619 ,
         \U1/aes_core/SB3/n2618 , \U1/aes_core/SB3/n2617 ,
         \U1/aes_core/SB3/n2616 , \U1/aes_core/SB3/n2615 ,
         \U1/aes_core/SB3/n2614 , \U1/aes_core/SB3/n2613 ,
         \U1/aes_core/SB3/n2612 , \U1/aes_core/SB3/n2611 ,
         \U1/aes_core/SB3/n2610 , \U1/aes_core/SB3/n2609 ,
         \U1/aes_core/SB3/n2608 , \U1/aes_core/SB3/n2607 ,
         \U1/aes_core/SB3/n2606 , \U1/aes_core/SB3/n2605 ,
         \U1/aes_core/SB3/n2604 , \U1/aes_core/SB3/n2603 ,
         \U1/aes_core/SB3/n2602 , \U1/aes_core/SB3/n2601 ,
         \U1/aes_core/SB3/n2600 , \U1/aes_core/SB3/n2599 ,
         \U1/aes_core/SB3/n2598 , \U1/aes_core/SB3/n2597 ,
         \U1/aes_core/SB3/n2596 , \U1/aes_core/SB3/n2595 ,
         \U1/aes_core/SB3/n2594 , \U1/aes_core/SB3/n2593 ,
         \U1/aes_core/SB3/n2592 , \U1/aes_core/SB3/n2591 ,
         \U1/aes_core/SB3/n2590 , \U1/aes_core/SB3/n2589 ,
         \U1/aes_core/SB3/n2588 , \U1/aes_core/SB3/n2587 ,
         \U1/aes_core/SB3/n2586 , \U1/aes_core/SB3/n2585 ,
         \U1/aes_core/SB3/n2584 , \U1/aes_core/SB3/n2583 ,
         \U1/aes_core/SB3/n2582 , \U1/aes_core/SB3/n2581 ,
         \U1/aes_core/SB3/n2580 , \U1/aes_core/SB3/n2579 ,
         \U1/aes_core/SB3/n2578 , \U1/aes_core/SB3/n2577 ,
         \U1/aes_core/SB3/n2576 , \U1/aes_core/SB3/n2575 ,
         \U1/aes_core/SB3/n2574 , \U1/aes_core/SB3/n2573 ,
         \U1/aes_core/SB3/n2572 , \U1/aes_core/SB3/n2571 ,
         \U1/aes_core/SB3/n2570 , \U1/aes_core/SB3/n2569 ,
         \U1/aes_core/SB3/n2568 , \U1/aes_core/SB3/n2567 ,
         \U1/aes_core/SB3/n2566 , \U1/aes_core/SB3/n2565 ,
         \U1/aes_core/SB3/n2564 , \U1/aes_core/SB3/n2563 ,
         \U1/aes_core/SB3/n2562 , \U1/aes_core/SB3/n2561 ,
         \U1/aes_core/SB3/n2560 , \U1/aes_core/SB3/n2559 ,
         \U1/aes_core/SB3/n2558 , \U1/aes_core/SB3/n2557 ,
         \U1/aes_core/SB3/n2556 , \U1/aes_core/SB3/n2555 ,
         \U1/aes_core/SB3/n2554 , \U1/aes_core/SB3/n2553 ,
         \U1/aes_core/SB3/n2552 , \U1/aes_core/SB3/n2551 ,
         \U1/aes_core/SB3/n2550 , \U1/aes_core/SB3/n2549 ,
         \U1/aes_core/SB3/n2548 , \U1/aes_core/SB3/n2547 ,
         \U1/aes_core/SB3/n2546 , \U1/aes_core/SB3/n2545 ,
         \U1/aes_core/SB3/n2544 , \U1/aes_core/SB3/n2543 ,
         \U1/aes_core/SB3/n2542 , \U1/aes_core/SB3/n2541 ,
         \U1/aes_core/SB3/n2540 , \U1/aes_core/SB3/n2539 ,
         \U1/aes_core/SB3/n2538 , \U1/aes_core/SB3/n2537 ,
         \U1/aes_core/SB3/n2536 , \U1/aes_core/SB3/n2535 ,
         \U1/aes_core/SB3/n2534 , \U1/aes_core/SB3/n2533 ,
         \U1/aes_core/SB3/n2532 , \U1/aes_core/SB3/n2531 ,
         \U1/aes_core/SB3/n2530 , \U1/aes_core/SB3/n2529 ,
         \U1/aes_core/SB3/n2528 , \U1/aes_core/SB3/n2527 ,
         \U1/aes_core/SB3/n2526 , \U1/aes_core/SB3/n2525 ,
         \U1/aes_core/SB3/n2524 , \U1/aes_core/SB3/n2523 ,
         \U1/aes_core/SB3/n2522 , \U1/aes_core/SB3/n2521 ,
         \U1/aes_core/SB3/n2520 , \U1/aes_core/SB3/n2519 ,
         \U1/aes_core/SB3/n2518 , \U1/aes_core/SB3/n2517 ,
         \U1/aes_core/SB3/n2516 , \U1/aes_core/SB3/n2515 ,
         \U1/aes_core/SB3/n2514 , \U1/aes_core/SB3/n2513 ,
         \U1/aes_core/SB3/n2512 , \U1/aes_core/SB3/n2511 ,
         \U1/aes_core/SB3/n2510 , \U1/aes_core/SB3/n2509 ,
         \U1/aes_core/SB3/n2508 , \U1/aes_core/SB3/n2507 ,
         \U1/aes_core/SB3/n2506 , \U1/aes_core/SB3/n2505 ,
         \U1/aes_core/SB3/n2504 , \U1/aes_core/SB3/n2503 ,
         \U1/aes_core/SB3/n2502 , \U1/aes_core/SB3/n2501 ,
         \U1/aes_core/SB3/n2500 , \U1/aes_core/SB3/n2499 ,
         \U1/aes_core/SB3/n2498 , \U1/aes_core/SB3/n2497 ,
         \U1/aes_core/SB3/n2496 , \U1/aes_core/SB3/n2495 ,
         \U1/aes_core/SB3/n2494 , \U1/aes_core/SB3/n2493 ,
         \U1/aes_core/SB3/n2492 , \U1/aes_core/SB3/n2491 ,
         \U1/aes_core/SB3/n2490 , \U1/aes_core/SB3/n2489 ,
         \U1/aes_core/SB3/n2488 , \U1/aes_core/SB3/n2487 ,
         \U1/aes_core/SB3/n2486 , \U1/aes_core/SB3/n2485 ,
         \U1/aes_core/SB3/n2484 , \U1/aes_core/SB3/n2483 ,
         \U1/aes_core/SB3/n2482 , \U1/aes_core/SB3/n2481 ,
         \U1/aes_core/SB3/n2480 , \U1/aes_core/SB3/n2479 ,
         \U1/aes_core/SB3/n2478 , \U1/aes_core/SB3/n2477 ,
         \U1/aes_core/SB3/n2476 , \U1/aes_core/SB3/n2475 ,
         \U1/aes_core/SB3/n2474 , \U1/aes_core/SB3/n2473 ,
         \U1/aes_core/SB3/n2472 , \U1/aes_core/SB3/n2471 ,
         \U1/aes_core/SB3/n2470 , \U1/aes_core/SB3/n2469 ,
         \U1/aes_core/SB3/n2468 , \U1/aes_core/SB3/n2467 ,
         \U1/aes_core/SB3/n2466 , \U1/aes_core/SB3/n2465 ,
         \U1/aes_core/SB3/n2464 , \U1/aes_core/SB3/n2463 ,
         \U1/aes_core/SB3/n2462 , \U1/aes_core/SB3/n2461 ,
         \U1/aes_core/SB3/n2460 , \U1/aes_core/SB3/n2459 ,
         \U1/aes_core/SB3/n2458 , \U1/aes_core/SB3/n2457 ,
         \U1/aes_core/SB3/n2456 , \U1/aes_core/SB3/n2455 ,
         \U1/aes_core/SB3/n2454 , \U1/aes_core/SB3/n2453 ,
         \U1/aes_core/SB3/n2452 , \U1/aes_core/SB3/n2451 ,
         \U1/aes_core/SB3/n2450 , \U1/aes_core/SB3/n2449 ,
         \U1/aes_core/SB3/n2448 , \U1/aes_core/SB3/n2447 ,
         \U1/aes_core/SB3/n2446 , \U1/aes_core/SB3/n2445 ,
         \U1/aes_core/SB3/n2444 , \U1/aes_core/SB3/n2443 ,
         \U1/aes_core/SB3/n2442 , \U1/aes_core/SB3/n2441 ,
         \U1/aes_core/SB3/n2440 , \U1/aes_core/SB3/n2439 ,
         \U1/aes_core/SB3/n2438 , \U1/aes_core/SB3/n2437 ,
         \U1/aes_core/SB3/n2436 , \U1/aes_core/SB3/n2435 ,
         \U1/aes_core/SB3/n2434 , \U1/aes_core/SB3/n2433 ,
         \U1/aes_core/SB3/n2432 , \U1/aes_core/SB3/n2431 ,
         \U1/aes_core/SB3/n2430 , \U1/aes_core/SB3/n2429 ,
         \U1/aes_core/SB3/n2428 , \U1/aes_core/SB3/n2427 ,
         \U1/aes_core/SB3/n2426 , \U1/aes_core/SB3/n2425 ,
         \U1/aes_core/SB3/n2424 , \U1/aes_core/SB3/n2423 ,
         \U1/aes_core/SB3/n2422 , \U1/aes_core/SB3/n2421 ,
         \U1/aes_core/SB3/n2420 , \U1/aes_core/SB3/n2419 ,
         \U1/aes_core/SB3/n2418 , \U1/aes_core/SB3/n2417 ,
         \U1/aes_core/SB3/n2416 , \U1/aes_core/SB3/n2415 ,
         \U1/aes_core/SB3/n2414 , \U1/aes_core/SB3/n2413 ,
         \U1/aes_core/SB3/n2412 , \U1/aes_core/SB3/n2411 ,
         \U1/aes_core/SB3/n2410 , \U1/aes_core/SB3/n2409 ,
         \U1/aes_core/SB3/n2408 , \U1/aes_core/SB3/n2407 ,
         \U1/aes_core/SB3/n2406 , \U1/aes_core/SB3/n2405 ,
         \U1/aes_core/SB3/n2404 , \U1/aes_core/SB3/n2403 ,
         \U1/aes_core/SB3/n2402 , \U1/aes_core/SB3/n2401 ,
         \U1/aes_core/SB3/n2400 , \U1/aes_core/SB3/n2399 ,
         \U1/aes_core/SB3/n2398 , \U1/aes_core/SB3/n2397 ,
         \U1/aes_core/SB3/n2396 , \U1/aes_core/SB3/n2395 ,
         \U1/aes_core/SB3/n2394 , \U1/aes_core/SB3/n2393 ,
         \U1/aes_core/SB3/n2392 , \U1/aes_core/SB3/n2391 ,
         \U1/aes_core/SB3/n2390 , \U1/aes_core/SB3/n2389 ,
         \U1/aes_core/SB3/n2388 , \U1/aes_core/SB3/n2387 ,
         \U1/aes_core/SB3/n2386 , \U1/aes_core/SB3/n2385 ,
         \U1/aes_core/SB3/n2384 , \U1/aes_core/SB3/n2383 ,
         \U1/aes_core/SB3/n2382 , \U1/aes_core/SB3/n2381 ,
         \U1/aes_core/SB3/n2380 , \U1/aes_core/SB3/n2379 ,
         \U1/aes_core/SB3/n2378 , \U1/aes_core/SB3/n2377 ,
         \U1/aes_core/SB3/n2376 , \U1/aes_core/SB3/n2375 ,
         \U1/aes_core/SB3/n2374 , \U1/aes_core/SB3/n2373 ,
         \U1/aes_core/SB3/n2372 , \U1/aes_core/SB3/n2371 ,
         \U1/aes_core/SB3/n2370 , \U1/aes_core/SB3/n2369 ,
         \U1/aes_core/SB3/n2368 , \U1/aes_core/SB3/n2367 ,
         \U1/aes_core/SB3/n2366 , \U1/aes_core/SB3/n2365 ,
         \U1/aes_core/SB3/n2364 , \U1/aes_core/SB3/n2363 ,
         \U1/aes_core/SB3/n2362 , \U1/aes_core/SB3/n2361 ,
         \U1/aes_core/SB3/n2360 , \U1/aes_core/SB3/n2359 ,
         \U1/aes_core/SB3/n2358 , \U1/aes_core/SB3/n2357 ,
         \U1/aes_core/SB3/n2356 , \U1/aes_core/SB3/n2355 ,
         \U1/aes_core/SB3/n2354 , \U1/aes_core/SB3/n2353 ,
         \U1/aes_core/SB3/n2352 , \U1/aes_core/SB3/n2351 ,
         \U1/aes_core/SB3/n2350 , \U1/aes_core/SB3/n2349 ,
         \U1/aes_core/SB3/n2348 , \U1/aes_core/SB3/n2347 ,
         \U1/aes_core/SB3/n2346 , \U1/aes_core/SB3/n2345 ,
         \U1/aes_core/SB3/n2344 , \U1/aes_core/SB3/n2343 ,
         \U1/aes_core/SB3/n2342 , \U1/aes_core/SB3/n2341 ,
         \U1/aes_core/SB3/n2340 , \U1/aes_core/SB3/n2339 ,
         \U1/aes_core/SB3/n2338 , \U1/aes_core/SB3/n2337 ,
         \U1/aes_core/SB3/n2336 , \U1/aes_core/SB3/n2335 ,
         \U1/aes_core/SB3/n2334 , \U1/aes_core/SB3/n2333 ,
         \U1/aes_core/SB3/n2332 , \U1/aes_core/SB3/n2331 ,
         \U1/aes_core/SB3/n2330 , \U1/aes_core/SB3/n2329 ,
         \U1/aes_core/SB3/n2328 , \U1/aes_core/SB3/n2327 ,
         \U1/aes_core/SB3/n2326 , \U1/aes_core/SB3/n2325 ,
         \U1/aes_core/SB3/n2324 , \U1/aes_core/SB3/n2323 ,
         \U1/aes_core/SB3/n2322 , \U1/aes_core/SB3/n2321 ,
         \U1/aes_core/SB3/n2320 , \U1/aes_core/SB3/n2319 ,
         \U1/aes_core/SB3/n2318 , \U1/aes_core/SB3/n2317 ,
         \U1/aes_core/SB3/n2316 , \U1/aes_core/SB3/n2315 ,
         \U1/aes_core/SB3/n2314 , \U1/aes_core/SB3/n2313 ,
         \U1/aes_core/SB3/n2312 , \U1/aes_core/SB3/n2311 ,
         \U1/aes_core/SB3/n2310 , \U1/aes_core/SB3/n2309 ,
         \U1/aes_core/SB3/n2308 , \U1/aes_core/SB3/n2307 ,
         \U1/aes_core/SB3/n2306 , \U1/aes_core/SB3/n2305 ,
         \U1/aes_core/SB3/n2304 , \U1/aes_core/SB3/n2303 ,
         \U1/aes_core/SB3/n2302 , \U1/aes_core/SB3/n2301 ,
         \U1/aes_core/SB3/n2300 , \U1/aes_core/SB3/n2299 ,
         \U1/aes_core/SB3/n2298 , \U1/aes_core/SB3/n2297 ,
         \U1/aes_core/SB3/n2296 , \U1/aes_core/SB3/n2295 ,
         \U1/aes_core/SB3/n2294 , \U1/aes_core/SB3/n2293 ,
         \U1/aes_core/SB3/n2292 , \U1/aes_core/SB3/n2291 ,
         \U1/aes_core/SB3/n2290 , \U1/aes_core/SB3/n2289 ,
         \U1/aes_core/SB3/n2288 , \U1/aes_core/SB3/n2287 ,
         \U1/aes_core/SB3/n2286 , \U1/aes_core/SB3/n2285 ,
         \U1/aes_core/SB3/n2284 , \U1/aes_core/SB3/n2283 ,
         \U1/aes_core/SB3/n2282 , \U1/aes_core/SB3/n2281 ,
         \U1/aes_core/SB3/n2280 , \U1/aes_core/SB3/n2279 ,
         \U1/aes_core/SB3/n2278 , \U1/aes_core/SB3/n2277 ,
         \U1/aes_core/SB3/n2276 , \U1/aes_core/SB3/n2275 ,
         \U1/aes_core/SB3/n2274 , \U1/aes_core/SB3/n2273 ,
         \U1/aes_core/SB3/n2272 , \U1/aes_core/SB3/n2271 ,
         \U1/aes_core/SB3/n2270 , \U1/aes_core/SB3/n2269 ,
         \U1/aes_core/SB3/n2268 , \U1/aes_core/SB3/n2267 ,
         \U1/aes_core/SB3/n2266 , \U1/aes_core/SB3/n2265 ,
         \U1/aes_core/SB3/n2264 , \U1/aes_core/SB3/n2263 ,
         \U1/aes_core/SB3/n2262 , \U1/aes_core/SB3/n2261 ,
         \U1/aes_core/SB3/n2260 , \U1/aes_core/SB3/n2259 ,
         \U1/aes_core/SB3/n2258 , \U1/aes_core/SB3/n2257 ,
         \U1/aes_core/SB3/n2256 , \U1/aes_core/SB3/n2255 ,
         \U1/aes_core/SB3/n2254 , \U1/aes_core/SB3/n2253 ,
         \U1/aes_core/SB3/n2252 , \U1/aes_core/SB3/n2251 ,
         \U1/aes_core/SB3/n2250 , \U1/aes_core/SB3/n2249 ,
         \U1/aes_core/SB3/n2248 , \U1/aes_core/SB3/n2247 ,
         \U1/aes_core/SB3/n2246 , \U1/aes_core/SB3/n2245 ,
         \U1/aes_core/SB3/n2244 , \U1/aes_core/SB3/n2243 ,
         \U1/aes_core/SB3/n2242 , \U1/aes_core/SB3/n2241 ,
         \U1/aes_core/SB3/n2240 , \U1/aes_core/SB3/n2239 ,
         \U1/aes_core/SB3/n2238 , \U1/aes_core/SB3/n2237 ,
         \U1/aes_core/SB3/n2236 , \U1/aes_core/SB3/n2235 ,
         \U1/aes_core/SB3/n2234 , \U1/aes_core/SB3/n2233 ,
         \U1/aes_core/SB3/n2232 , \U1/aes_core/SB3/n2231 ,
         \U1/aes_core/SB3/n2230 , \U1/aes_core/SB3/n2229 ,
         \U1/aes_core/SB3/n2228 , \U1/aes_core/SB3/n2227 ,
         \U1/aes_core/SB3/n2226 , \U1/aes_core/SB3/n2225 ,
         \U1/aes_core/SB3/n2224 , \U1/aes_core/SB3/n2223 ,
         \U1/aes_core/SB3/n2222 , \U1/aes_core/SB3/n2221 ,
         \U1/aes_core/SB3/n2220 , \U1/aes_core/SB3/n2219 ,
         \U1/aes_core/SB3/n2218 , \U1/aes_core/SB3/n2217 ,
         \U1/aes_core/SB3/n2216 , \U1/aes_core/SB3/n2215 ,
         \U1/aes_core/SB3/n2214 , \U1/aes_core/SB3/n2213 ,
         \U1/aes_core/SB3/n2212 , \U1/aes_core/SB3/n2211 ,
         \U1/aes_core/SB3/n2210 , \U1/aes_core/SB3/n2209 ,
         \U1/aes_core/SB3/n2208 , \U1/aes_core/SB3/n2207 ,
         \U1/aes_core/SB3/n2206 , \U1/aes_core/SB3/n2205 ,
         \U1/aes_core/SB3/n2204 , \U1/aes_core/SB3/n2203 ,
         \U1/aes_core/SB3/n2202 , \U1/aes_core/SB3/n2201 ,
         \U1/aes_core/SB3/n2200 , \U1/aes_core/SB3/n2199 ,
         \U1/aes_core/SB3/n2198 , \U1/aes_core/SB3/n2197 ,
         \U1/aes_core/SB3/n2196 , \U1/aes_core/SB3/n2195 ,
         \U1/aes_core/SB3/n2194 , \U1/aes_core/SB3/n2193 ,
         \U1/aes_core/SB3/n2192 , \U1/aes_core/SB3/n2191 ,
         \U1/aes_core/SB3/n2190 , \U1/aes_core/SB3/n2189 ,
         \U1/aes_core/SB3/n2188 , \U1/aes_core/SB3/n2187 ,
         \U1/aes_core/SB3/n2186 , \U1/aes_core/SB3/n2185 ,
         \U1/aes_core/SB3/n2184 , \U1/aes_core/SB3/n2183 ,
         \U1/aes_core/SB3/n2182 , \U1/aes_core/SB3/n2181 ,
         \U1/aes_core/SB3/n2180 , \U1/aes_core/SB3/n2179 ,
         \U1/aes_core/SB3/n2178 , \U1/aes_core/SB3/n2177 ,
         \U1/aes_core/SB3/n2176 , \U1/aes_core/SB3/n2175 ,
         \U1/aes_core/SB3/n2174 , \U1/aes_core/SB3/n2173 ,
         \U1/aes_core/SB3/n2172 , \U1/aes_core/SB3/n2171 ,
         \U1/aes_core/SB3/n2170 , \U1/aes_core/SB3/n2169 ,
         \U1/aes_core/SB3/n2168 , \U1/aes_core/SB3/n2167 ,
         \U1/aes_core/SB3/n2166 , \U1/aes_core/SB3/n2165 ,
         \U1/aes_core/SB3/n2164 , \U1/aes_core/SB3/n2163 ,
         \U1/aes_core/SB3/n2162 , \U1/aes_core/SB3/n2161 ,
         \U1/aes_core/SB3/n2160 , \U1/aes_core/SB3/n2159 ,
         \U1/aes_core/SB3/n2158 , \U1/aes_core/SB3/n2157 ,
         \U1/aes_core/SB3/n2156 , \U1/aes_core/SB3/n2155 ,
         \U1/aes_core/SB3/n2154 , \U1/aes_core/SB3/n2153 ,
         \U1/aes_core/SB3/n2152 , \U1/aes_core/SB3/n2151 ,
         \U1/aes_core/SB3/n2150 , \U1/aes_core/SB3/n2149 ,
         \U1/aes_core/SB3/n2148 , \U1/aes_core/SB3/n2147 ,
         \U1/aes_core/SB3/n2146 , \U1/aes_core/SB3/n2145 ,
         \U1/aes_core/SB3/n2144 , \U1/aes_core/SB3/n2143 ,
         \U1/aes_core/SB3/n2142 , \U1/aes_core/SB3/n2141 ,
         \U1/aes_core/SB3/n2140 , \U1/aes_core/SB3/n2139 ,
         \U1/aes_core/SB3/n2138 , \U1/aes_core/SB3/n2137 ,
         \U1/aes_core/SB3/n2136 , \U1/aes_core/SB3/n2135 ,
         \U1/aes_core/SB3/n2134 , \U1/aes_core/SB3/n2133 ,
         \U1/aes_core/SB3/n2132 , \U1/aes_core/SB3/n2131 ,
         \U1/aes_core/SB3/n2130 , \U1/aes_core/SB3/n2129 ,
         \U1/aes_core/SB3/n2128 , \U1/aes_core/SB3/n2127 ,
         \U1/aes_core/SB3/n2126 , \U1/aes_core/SB3/n2125 ,
         \U1/aes_core/SB3/n2124 , \U1/aes_core/SB3/n2123 ,
         \U1/aes_core/SB3/n2122 , \U1/aes_core/SB3/n2121 ,
         \U1/aes_core/SB3/n2120 , \U1/aes_core/SB3/n2119 ,
         \U1/aes_core/SB3/n2118 , \U1/aes_core/SB3/n2117 ,
         \U1/aes_core/SB3/n2116 , \U1/aes_core/SB3/n2115 ,
         \U1/aes_core/SB3/n2114 , \U1/aes_core/SB3/n2113 ,
         \U1/aes_core/SB3/n2112 , \U1/aes_core/SB3/n2111 ,
         \U1/aes_core/SB3/n2110 , \U1/aes_core/SB3/n2109 ,
         \U1/aes_core/SB3/n2108 , \U1/aes_core/SB3/n2107 ,
         \U1/aes_core/SB3/n2106 , \U1/aes_core/SB3/n2105 ,
         \U1/aes_core/SB3/n2104 , \U1/aes_core/SB3/n2103 ,
         \U1/aes_core/SB3/n2102 , \U1/aes_core/SB3/n2101 ,
         \U1/aes_core/SB3/n2100 , \U1/aes_core/SB3/n2099 ,
         \U1/aes_core/SB3/n2098 , \U1/aes_core/SB3/n2097 ,
         \U1/aes_core/SB3/n2096 , \U1/aes_core/SB3/n2095 ,
         \U1/aes_core/SB3/n2094 , \U1/aes_core/SB3/n2093 ,
         \U1/aes_core/SB3/n2092 , \U1/aes_core/SB3/n2091 ,
         \U1/aes_core/SB3/n2090 , \U1/aes_core/SB3/n2089 ,
         \U1/aes_core/SB3/n2088 , \U1/aes_core/SB3/n2087 ,
         \U1/aes_core/SB3/n2086 , \U1/aes_core/SB3/n2085 ,
         \U1/aes_core/SB3/n2084 , \U1/aes_core/SB3/n2083 ,
         \U1/aes_core/SB3/n2082 , \U1/aes_core/SB3/n2081 ,
         \U1/aes_core/SB3/n2080 , \U1/aes_core/SB3/n2079 ,
         \U1/aes_core/SB3/n2078 , \U1/aes_core/SB3/n2077 ,
         \U1/aes_core/SB3/n2076 , \U1/aes_core/SB3/n2075 ,
         \U1/aes_core/SB3/n2074 , \U1/aes_core/SB3/n2073 ,
         \U1/aes_core/SB3/n2072 , \U1/aes_core/SB3/n2071 ,
         \U1/aes_core/SB3/n2070 , \U1/aes_core/SB3/n2069 ,
         \U1/aes_core/SB3/n2068 , \U1/aes_core/SB3/n2067 ,
         \U1/aes_core/SB3/n2066 , \U1/aes_core/SB3/n2065 ,
         \U1/aes_core/SB3/n2064 , \U1/aes_core/SB3/n2063 ,
         \U1/aes_core/SB3/n2062 , \U1/aes_core/SB3/n2061 ,
         \U1/aes_core/SB3/n2060 , \U1/aes_core/SB3/n2059 ,
         \U1/aes_core/SB3/n2058 , \U1/aes_core/SB3/n2057 ,
         \U1/aes_core/SB3/n2056 , \U1/aes_core/SB3/n2055 ,
         \U1/aes_core/SB3/n2054 , \U1/aes_core/SB3/n2053 ,
         \U1/aes_core/SB3/n2052 , \U1/aes_core/SB3/n2051 ,
         \U1/aes_core/SB3/n2050 , \U1/aes_core/SB3/n2049 ,
         \U1/aes_core/SB3/n2048 , \U1/aes_core/SB3/n2047 ,
         \U1/aes_core/SB3/n2046 , \U1/aes_core/SB3/n2045 ,
         \U1/aes_core/SB3/n2044 , \U1/aes_core/SB3/n2043 ,
         \U1/aes_core/SB3/n2042 , \U1/aes_core/SB3/n2041 ,
         \U1/aes_core/SB3/n2040 , \U1/aes_core/SB3/n2039 ,
         \U1/aes_core/SB3/n2038 , \U1/aes_core/SB3/n2037 ,
         \U1/aes_core/SB3/n2036 , \U1/aes_core/SB3/n2035 ,
         \U1/aes_core/SB3/n2034 , \U1/aes_core/SB3/n2033 ,
         \U1/aes_core/SB3/n2032 , \U1/aes_core/SB3/n2031 ,
         \U1/aes_core/SB3/n2030 , \U1/aes_core/SB3/n2029 ,
         \U1/aes_core/SB3/n2028 , \U1/aes_core/SB3/n2027 ,
         \U1/aes_core/SB3/n2026 , \U1/aes_core/SB3/n2025 ,
         \U1/aes_core/SB3/n2024 , \U1/aes_core/SB3/n2023 ,
         \U1/aes_core/SB3/n2022 , \U1/aes_core/SB3/n2021 ,
         \U1/aes_core/SB3/n2020 , \U1/aes_core/SB3/n2019 ,
         \U1/aes_core/SB3/n2018 , \U1/aes_core/SB3/n2017 ,
         \U1/aes_core/SB3/n2016 , \U1/aes_core/SB3/n2015 ,
         \U1/aes_core/SB3/n2014 , \U1/aes_core/SB3/n2013 ,
         \U1/aes_core/SB3/n2012 , \U1/aes_core/SB3/n2011 ,
         \U1/aes_core/SB3/n2010 , \U1/aes_core/SB3/n2009 ,
         \U1/aes_core/SB3/n2008 , \U1/aes_core/SB3/n2007 ,
         \U1/aes_core/SB3/n2006 , \U1/aes_core/SB3/n2005 ,
         \U1/aes_core/SB3/n2004 , \U1/aes_core/SB3/n2003 ,
         \U1/aes_core/SB3/n2002 , \U1/aes_core/SB3/n2001 ,
         \U1/aes_core/SB3/n2000 , \U1/aes_core/SB3/n1999 ,
         \U1/aes_core/SB3/n1998 , \U1/aes_core/SB3/n1997 ,
         \U1/aes_core/SB3/n1996 , \U1/aes_core/SB3/n1995 ,
         \U1/aes_core/SB3/n1994 , \U1/aes_core/SB3/n1993 ,
         \U1/aes_core/SB3/n1992 , \U1/aes_core/SB3/n1991 ,
         \U1/aes_core/SB3/n1990 , \U1/aes_core/SB3/n1989 ,
         \U1/aes_core/SB3/n1988 , \U1/aes_core/SB3/n1987 ,
         \U1/aes_core/SB3/n1986 , \U1/aes_core/SB3/n1985 ,
         \U1/aes_core/SB3/n1984 , \U1/aes_core/SB3/n1983 ,
         \U1/aes_core/SB3/n1982 , \U1/aes_core/SB3/n1981 ,
         \U1/aes_core/SB3/n1980 , \U1/aes_core/SB3/n1979 ,
         \U1/aes_core/SB3/n1978 , \U1/aes_core/SB3/n1977 ,
         \U1/aes_core/SB3/n1976 , \U1/aes_core/SB3/n1975 ,
         \U1/aes_core/SB3/n1974 , \U1/aes_core/SB3/n1973 ,
         \U1/aes_core/SB3/n1972 , \U1/aes_core/SB3/n1971 ,
         \U1/aes_core/SB3/n1970 , \U1/aes_core/SB3/n1969 ,
         \U1/aes_core/SB3/n1968 , \U1/aes_core/SB3/n1967 ,
         \U1/aes_core/SB3/n1966 , \U1/aes_core/SB3/n1965 ,
         \U1/aes_core/SB3/n1964 , \U1/aes_core/SB3/n1963 ,
         \U1/aes_core/SB3/n1962 , \U1/aes_core/SB3/n1961 ,
         \U1/aes_core/SB3/n1960 , \U1/aes_core/SB3/n1959 ,
         \U1/aes_core/SB3/n1958 , \U1/aes_core/SB3/n1957 ,
         \U1/aes_core/SB3/n1956 , \U1/aes_core/SB3/n1955 ,
         \U1/aes_core/SB3/n1954 , \U1/aes_core/SB3/n1953 ,
         \U1/aes_core/SB3/n1952 , \U1/aes_core/SB3/n1951 ,
         \U1/aes_core/SB3/n1950 , \U1/aes_core/SB3/n1949 ,
         \U1/aes_core/SB3/n1948 , \U1/aes_core/SB3/n1947 ,
         \U1/aes_core/SB3/n1946 , \U1/aes_core/SB3/n1945 ,
         \U1/aes_core/SB3/n1944 , \U1/aes_core/SB3/n1943 ,
         \U1/aes_core/SB3/n1942 , \U1/aes_core/SB3/n1941 ,
         \U1/aes_core/SB3/n1940 , \U1/aes_core/SB3/n1939 ,
         \U1/aes_core/SB3/n1938 , \U1/aes_core/SB3/n1937 ,
         \U1/aes_core/SB3/n1936 , \U1/aes_core/SB3/n1935 ,
         \U1/aes_core/SB3/n1934 , \U1/aes_core/SB3/n1933 ,
         \U1/aes_core/SB3/n1932 , \U1/aes_core/SB3/n1931 ,
         \U1/aes_core/SB3/n1930 , \U1/aes_core/SB3/n1929 ,
         \U1/aes_core/SB3/n1928 , \U1/aes_core/SB3/n1927 ,
         \U1/aes_core/SB3/n1926 , \U1/aes_core/SB3/n1925 ,
         \U1/aes_core/SB3/n1924 , \U1/aes_core/SB3/n1923 ,
         \U1/aes_core/SB3/n1922 , \U1/aes_core/SB3/n1921 ,
         \U1/aes_core/SB3/n1920 , \U1/aes_core/SB3/n1919 ,
         \U1/aes_core/SB3/n1918 , \U1/aes_core/SB3/n1917 ,
         \U1/aes_core/SB3/n1916 , \U1/aes_core/SB3/n1915 ,
         \U1/aes_core/SB3/n1914 , \U1/aes_core/SB3/n1913 ,
         \U1/aes_core/SB3/n1912 , \U1/aes_core/SB3/n1911 ,
         \U1/aes_core/SB3/n1910 , \U1/aes_core/SB3/n1909 ,
         \U1/aes_core/SB3/n1908 , \U1/aes_core/SB3/n1907 ,
         \U1/aes_core/SB3/n1906 , \U1/aes_core/SB3/n1905 ,
         \U1/aes_core/SB3/n1904 , \U1/aes_core/SB3/n1903 ,
         \U1/aes_core/SB3/n1902 , \U1/aes_core/SB3/n1901 ,
         \U1/aes_core/SB3/n1900 , \U1/aes_core/SB3/n1899 ,
         \U1/aes_core/SB3/n1898 , \U1/aes_core/SB3/n1897 ,
         \U1/aes_core/SB3/n1896 , \U1/aes_core/SB3/n1895 ,
         \U1/aes_core/SB3/n1894 , \U1/aes_core/SB3/n1893 ,
         \U1/aes_core/SB3/n1892 , \U1/aes_core/SB3/n1891 ,
         \U1/aes_core/SB3/n1890 , \U1/aes_core/SB3/n1889 ,
         \U1/aes_core/SB3/n1888 , \U1/aes_core/SB3/n1887 ,
         \U1/aes_core/SB3/n1886 , \U1/aes_core/SB3/n1885 ,
         \U1/aes_core/SB3/n1884 , \U1/aes_core/SB3/n1883 ,
         \U1/aes_core/SB3/n1882 , \U1/aes_core/SB3/n1881 ,
         \U1/aes_core/SB3/n1880 , \U1/aes_core/SB3/n1879 ,
         \U1/aes_core/SB3/n1878 , \U1/aes_core/SB3/n1877 ,
         \U1/aes_core/SB3/n1876 , \U1/aes_core/SB3/n1875 ,
         \U1/aes_core/SB3/n1874 , \U1/aes_core/SB3/n1873 ,
         \U1/aes_core/SB3/n1872 , \U1/aes_core/SB3/n1871 ,
         \U1/aes_core/SB3/n1870 , \U1/aes_core/SB3/n1869 ,
         \U1/aes_core/SB3/n1868 , \U1/aes_core/SB3/n1867 ,
         \U1/aes_core/SB3/n1866 , \U1/aes_core/SB3/n1865 ,
         \U1/aes_core/SB3/n1864 , \U1/aes_core/SB3/n1863 ,
         \U1/aes_core/SB3/n1862 , \U1/aes_core/SB3/n1861 ,
         \U1/aes_core/SB3/n1860 , \U1/aes_core/SB3/n1859 ,
         \U1/aes_core/SB3/n1858 , \U1/aes_core/SB3/n1857 ,
         \U1/aes_core/SB3/n1856 , \U1/aes_core/SB3/n1855 ,
         \U1/aes_core/SB3/n1854 , \U1/aes_core/SB3/n1853 ,
         \U1/aes_core/SB3/n1852 , \U1/aes_core/SB3/n1851 ,
         \U1/aes_core/SB3/n1850 , \U1/aes_core/SB3/n1849 ,
         \U1/aes_core/SB3/n1848 , \U1/aes_core/SB3/n1847 ,
         \U1/aes_core/SB3/n1846 , \U1/aes_core/SB3/n1845 ,
         \U1/aes_core/SB3/n1844 , \U1/aes_core/SB3/n1843 ,
         \U1/aes_core/SB3/n1842 , \U1/aes_core/SB3/n1841 ,
         \U1/aes_core/SB3/n1840 , \U1/aes_core/SB3/n1839 ,
         \U1/aes_core/SB3/n1838 , \U1/aes_core/SB3/n1837 ,
         \U1/aes_core/SB3/n1836 , \U1/aes_core/SB3/n1835 ,
         \U1/aes_core/SB3/n1834 , \U1/aes_core/SB3/n1833 ,
         \U1/aes_core/SB3/n1832 , \U1/aes_core/SB3/n1831 ,
         \U1/aes_core/SB3/n1830 , \U1/aes_core/SB3/n1829 ,
         \U1/aes_core/SB3/n1828 , \U1/aes_core/SB3/n1827 ,
         \U1/aes_core/SB3/n1826 , \U1/aes_core/SB3/n1825 ,
         \U1/aes_core/SB3/n1824 , \U1/aes_core/SB3/n1823 ,
         \U1/aes_core/SB3/n1822 , \U1/aes_core/SB3/n1821 ,
         \U1/aes_core/SB3/n1820 , \U1/aes_core/SB3/n1819 ,
         \U1/aes_core/SB3/n1818 , \U1/aes_core/SB3/n1817 ,
         \U1/aes_core/SB3/n1816 , \U1/aes_core/SB3/n1815 ,
         \U1/aes_core/SB3/n1814 , \U1/aes_core/SB3/n1813 ,
         \U1/aes_core/SB3/n1812 , \U1/aes_core/SB3/n1811 ,
         \U1/aes_core/SB3/n1810 , \U1/aes_core/SB3/n1809 ,
         \U1/aes_core/SB3/n1808 , \U1/aes_core/SB3/n1807 ,
         \U1/aes_core/SB3/n1806 , \U1/aes_core/SB3/n1805 ,
         \U1/aes_core/SB3/n1804 , \U1/aes_core/SB3/n1803 ,
         \U1/aes_core/SB3/n1802 , \U1/aes_core/SB3/n1801 ,
         \U1/aes_core/SB3/n1800 , \U1/aes_core/SB3/n1799 ,
         \U1/aes_core/SB3/n1798 , \U1/aes_core/SB3/n1797 ,
         \U1/aes_core/SB3/n1796 , \U1/aes_core/SB3/n1795 ,
         \U1/aes_core/SB3/n1794 , \U1/aes_core/SB3/n1793 ,
         \U1/aes_core/SB3/n1792 , \U1/aes_core/SB3/n1791 ,
         \U1/aes_core/SB3/n1790 , \U1/aes_core/SB3/n1789 ,
         \U1/aes_core/SB3/n1788 , \U1/aes_core/SB3/n1787 ,
         \U1/aes_core/SB3/n1786 , \U1/aes_core/SB3/n1785 ,
         \U1/aes_core/SB3/n1784 , \U1/aes_core/SB3/n1783 ,
         \U1/aes_core/SB3/n1782 , \U1/aes_core/SB3/n1781 ,
         \U1/aes_core/SB3/n1780 , \U1/aes_core/SB3/n1779 ,
         \U1/aes_core/SB3/n1778 , \U1/aes_core/SB3/n1777 ,
         \U1/aes_core/SB3/n1776 , \U1/aes_core/SB3/n1775 ,
         \U1/aes_core/SB3/n1774 , \U1/aes_core/SB3/n1773 ,
         \U1/aes_core/SB3/n1772 , \U1/aes_core/SB3/n1771 ,
         \U1/aes_core/SB3/n1770 , \U1/aes_core/SB3/n1769 ,
         \U1/aes_core/SB3/n1768 , \U1/aes_core/SB3/n1767 ,
         \U1/aes_core/SB3/n1766 , \U1/aes_core/SB3/n1765 ,
         \U1/aes_core/SB3/n1764 , \U1/aes_core/SB3/n1763 ,
         \U1/aes_core/SB3/n1762 , \U1/aes_core/SB3/n1761 ,
         \U1/aes_core/SB3/n1760 , \U1/aes_core/SB3/n1759 ,
         \U1/aes_core/SB3/n1758 , \U1/aes_core/SB3/n1757 ,
         \U1/aes_core/SB3/n1756 , \U1/aes_core/SB3/n1755 ,
         \U1/aes_core/SB3/n1754 , \U1/aes_core/SB3/n1753 ,
         \U1/aes_core/SB3/n1752 , \U1/aes_core/SB3/n1751 ,
         \U1/aes_core/SB3/n1750 , \U1/aes_core/SB3/n1749 ,
         \U1/aes_core/SB3/n1748 , \U1/aes_core/SB3/n1747 ,
         \U1/aes_core/SB3/n1746 , \U1/aes_core/SB3/n1745 ,
         \U1/aes_core/SB3/n1744 , \U1/aes_core/SB3/n1743 ,
         \U1/aes_core/SB3/n1742 , \U1/aes_core/SB3/n1741 ,
         \U1/aes_core/SB3/n1740 , \U1/aes_core/SB3/n1739 ,
         \U1/aes_core/SB3/n1738 , \U1/aes_core/SB3/n1737 ,
         \U1/aes_core/SB3/n1736 , \U1/aes_core/SB3/n1735 ,
         \U1/aes_core/SB3/n1734 , \U1/aes_core/SB3/n1733 ,
         \U1/aes_core/SB3/n1732 , \U1/aes_core/SB3/n1731 ,
         \U1/aes_core/SB3/n1730 , \U1/aes_core/SB3/n1729 ,
         \U1/aes_core/SB3/n1728 , \U1/aes_core/SB3/n1727 ,
         \U1/aes_core/SB3/n1726 , \U1/aes_core/SB3/n1725 ,
         \U1/aes_core/SB3/n1724 , \U1/aes_core/SB3/n1723 ,
         \U1/aes_core/SB3/n1722 , \U1/aes_core/SB3/n1721 ,
         \U1/aes_core/SB3/n1720 , \U1/aes_core/SB3/n1719 ,
         \U1/aes_core/SB3/n1718 , \U1/aes_core/SB3/n1717 ,
         \U1/aes_core/SB3/n1716 , \U1/aes_core/SB3/n1715 ,
         \U1/aes_core/SB3/n1714 , \U1/aes_core/SB3/n1713 ,
         \U1/aes_core/SB3/n1712 , \U1/aes_core/SB3/n1711 ,
         \U1/aes_core/SB3/n1710 , \U1/aes_core/SB3/n1709 ,
         \U1/aes_core/SB3/n1708 , \U1/aes_core/SB3/n1707 ,
         \U1/aes_core/SB3/n1706 , \U1/aes_core/SB3/n1705 ,
         \U1/aes_core/SB3/n1704 , \U1/aes_core/SB3/n1703 ,
         \U1/aes_core/SB3/n1702 , \U1/aes_core/SB3/n1701 ,
         \U1/aes_core/SB3/n1700 , \U1/aes_core/SB3/n1699 ,
         \U1/aes_core/SB3/n1698 , \U1/aes_core/SB3/n1697 ,
         \U1/aes_core/SB3/n1696 , \U1/aes_core/SB3/n1695 ,
         \U1/aes_core/SB3/n1694 , \U1/aes_core/SB3/n1693 ,
         \U1/aes_core/SB3/n1692 , \U1/aes_core/SB3/n1691 ,
         \U1/aes_core/SB3/n1690 , \U1/aes_core/SB3/n1689 ,
         \U1/aes_core/SB3/n1688 , \U1/aes_core/SB3/n1687 ,
         \U1/aes_core/SB3/n1686 , \U1/aes_core/SB3/n1685 ,
         \U1/aes_core/SB3/n1684 , \U1/aes_core/SB3/n1683 ,
         \U1/aes_core/SB3/n1682 , \U1/aes_core/SB3/n1621 ,
         \U1/aes_core/SB3/n1218 , \U1/aes_core/SB3/n1203 ,
         \U1/aes_core/SB3/n1158 , \U1/aes_core/SB3/n1030 ,
         \U1/aes_core/SB3/n767 , \U1/aes_core/SB3/n752 ,
         \U1/aes_core/SB3/n707 , \U1/aes_core/SB3/n385 , \U1/aes_core/MC0/n80 ,
         \U1/aes_core/MC0/n79 , \U1/aes_core/MC0/n78 , \U1/aes_core/MC0/n77 ,
         \U1/aes_core/MC0/n76 , \U1/aes_core/MC0/n75 , \U1/aes_core/MC0/n74 ,
         \U1/aes_core/MC0/n73 , \U1/aes_core/MC0/n72 , \U1/aes_core/MC0/n71 ,
         \U1/aes_core/MC0/n70 , \U1/aes_core/MC0/n69 , \U1/aes_core/MC0/n68 ,
         \U1/aes_core/MC0/n67 , \U1/aes_core/MC0/n66 , \U1/aes_core/MC0/n65 ,
         \U1/aes_core/MC0/n64 , \U1/aes_core/MC0/n63 , \U1/aes_core/MC0/n62 ,
         \U1/aes_core/MC0/n61 , \U1/aes_core/MC0/n60 , \U1/aes_core/MC0/n59 ,
         \U1/aes_core/MC0/n58 , \U1/aes_core/MC0/n57 , \U1/aes_core/MC0/n56 ,
         \U1/aes_core/MC0/n55 , \U1/aes_core/MC0/n54 , \U1/aes_core/MC0/n53 ,
         \U1/aes_core/MC0/n52 , \U1/aes_core/MC0/n51 , \U1/aes_core/MC0/n50 ,
         \U1/aes_core/MC0/n49 , \U1/aes_core/MC0/n48 , \U1/aes_core/MC0/n47 ,
         \U1/aes_core/MC0/n46 , \U1/aes_core/MC0/n45 , \U1/aes_core/MC0/n44 ,
         \U1/aes_core/MC0/n43 , \U1/aes_core/MC0/n42 , \U1/aes_core/MC0/n41 ,
         \U1/aes_core/MC0/n40 , \U1/aes_core/MC0/n39 , \U1/aes_core/MC0/n38 ,
         \U1/aes_core/MC0/n36 , \U1/aes_core/MC0/n35 , \U1/aes_core/MC0/n33 ,
         \U1/aes_core/MC0/n32 , \U1/aes_core/MC0/n31 , \U1/aes_core/MC0/n30 ,
         \U1/aes_core/MC0/n29 , \U1/aes_core/MC0/n28 , \U1/aes_core/MC0/n27 ,
         \U1/aes_core/MC0/n26 , \U1/aes_core/MC0/n25 , \U1/aes_core/MC0/n24 ,
         \U1/aes_core/MC0/n23 , \U1/aes_core/MC0/n22 , \U1/aes_core/MC0/n21 ,
         \U1/aes_core/MC0/n20 , \U1/aes_core/MC0/n19 , \U1/aes_core/MC0/n18 ,
         \U1/aes_core/MC0/n17 , \U1/aes_core/MC0/n16 , \U1/aes_core/MC0/n15 ,
         \U1/aes_core/MC0/n14 , \U1/aes_core/MC0/n13 , \U1/aes_core/MC0/n12 ,
         \U1/aes_core/MC0/n11 , \U1/aes_core/MC0/n10 , \U1/aes_core/MC0/n9 ,
         \U1/aes_core/MC0/n8 , \U1/aes_core/MC0/n7 , \U1/aes_core/MC0/n6 ,
         \U1/aes_core/MC0/n5 , \U1/aes_core/MC0/n4 , \U1/aes_core/MC0/n3 ,
         \U1/aes_core/MC0/n2 , \U1/aes_core/MC1/n151 , \U1/aes_core/MC1/n150 ,
         \U1/aes_core/MC1/n149 , \U1/aes_core/MC1/n148 ,
         \U1/aes_core/MC1/n147 , \U1/aes_core/MC1/n146 ,
         \U1/aes_core/MC1/n145 , \U1/aes_core/MC1/n144 ,
         \U1/aes_core/MC1/n143 , \U1/aes_core/MC1/n142 ,
         \U1/aes_core/MC1/n141 , \U1/aes_core/MC1/n140 ,
         \U1/aes_core/MC1/n139 , \U1/aes_core/MC1/n138 ,
         \U1/aes_core/MC1/n137 , \U1/aes_core/MC1/n136 ,
         \U1/aes_core/MC1/n135 , \U1/aes_core/MC1/n134 ,
         \U1/aes_core/MC1/n133 , \U1/aes_core/MC1/n132 ,
         \U1/aes_core/MC1/n131 , \U1/aes_core/MC1/n130 ,
         \U1/aes_core/MC1/n129 , \U1/aes_core/MC1/n128 ,
         \U1/aes_core/MC1/n127 , \U1/aes_core/MC1/n126 ,
         \U1/aes_core/MC1/n125 , \U1/aes_core/MC1/n124 ,
         \U1/aes_core/MC1/n123 , \U1/aes_core/MC1/n122 ,
         \U1/aes_core/MC1/n121 , \U1/aes_core/MC1/n120 ,
         \U1/aes_core/MC1/n119 , \U1/aes_core/MC1/n118 ,
         \U1/aes_core/MC1/n117 , \U1/aes_core/MC1/n116 ,
         \U1/aes_core/MC1/n115 , \U1/aes_core/MC1/n114 ,
         \U1/aes_core/MC1/n113 , \U1/aes_core/MC1/n112 ,
         \U1/aes_core/MC1/n111 , \U1/aes_core/MC1/n110 ,
         \U1/aes_core/MC1/n109 , \U1/aes_core/MC1/n108 ,
         \U1/aes_core/MC1/n107 , \U1/aes_core/MC1/n106 ,
         \U1/aes_core/MC1/n105 , \U1/aes_core/MC1/n104 ,
         \U1/aes_core/MC1/n103 , \U1/aes_core/MC1/n102 ,
         \U1/aes_core/MC1/n101 , \U1/aes_core/MC1/n100 , \U1/aes_core/MC1/n99 ,
         \U1/aes_core/MC1/n98 , \U1/aes_core/MC1/n97 , \U1/aes_core/MC1/n96 ,
         \U1/aes_core/MC1/n95 , \U1/aes_core/MC1/n94 , \U1/aes_core/MC1/n93 ,
         \U1/aes_core/MC1/n92 , \U1/aes_core/MC1/n91 , \U1/aes_core/MC1/n90 ,
         \U1/aes_core/MC1/n89 , \U1/aes_core/MC1/n88 , \U1/aes_core/MC1/n87 ,
         \U1/aes_core/MC1/n86 , \U1/aes_core/MC1/n85 , \U1/aes_core/MC1/n84 ,
         \U1/aes_core/MC1/n83 , \U1/aes_core/MC1/n82 , \U1/aes_core/MC1/n81 ,
         \U1/aes_core/MC1/n80 , \U1/aes_core/MC1/n79 , \U1/aes_core/MC1/n78 ,
         \U1/aes_core/MC1/n37 , \U1/aes_core/MC1/n34 , \U1/aes_core/MC1/n1 ,
         \U1/aes_core/MC2/n151 , \U1/aes_core/MC2/n150 ,
         \U1/aes_core/MC2/n149 , \U1/aes_core/MC2/n148 ,
         \U1/aes_core/MC2/n147 , \U1/aes_core/MC2/n146 ,
         \U1/aes_core/MC2/n145 , \U1/aes_core/MC2/n144 ,
         \U1/aes_core/MC2/n143 , \U1/aes_core/MC2/n142 ,
         \U1/aes_core/MC2/n141 , \U1/aes_core/MC2/n140 ,
         \U1/aes_core/MC2/n139 , \U1/aes_core/MC2/n138 ,
         \U1/aes_core/MC2/n137 , \U1/aes_core/MC2/n136 ,
         \U1/aes_core/MC2/n135 , \U1/aes_core/MC2/n134 ,
         \U1/aes_core/MC2/n133 , \U1/aes_core/MC2/n132 ,
         \U1/aes_core/MC2/n131 , \U1/aes_core/MC2/n130 ,
         \U1/aes_core/MC2/n129 , \U1/aes_core/MC2/n128 ,
         \U1/aes_core/MC2/n127 , \U1/aes_core/MC2/n126 ,
         \U1/aes_core/MC2/n125 , \U1/aes_core/MC2/n124 ,
         \U1/aes_core/MC2/n123 , \U1/aes_core/MC2/n122 ,
         \U1/aes_core/MC2/n121 , \U1/aes_core/MC2/n120 ,
         \U1/aes_core/MC2/n119 , \U1/aes_core/MC2/n118 ,
         \U1/aes_core/MC2/n117 , \U1/aes_core/MC2/n116 ,
         \U1/aes_core/MC2/n115 , \U1/aes_core/MC2/n114 ,
         \U1/aes_core/MC2/n113 , \U1/aes_core/MC2/n112 ,
         \U1/aes_core/MC2/n111 , \U1/aes_core/MC2/n110 ,
         \U1/aes_core/MC2/n109 , \U1/aes_core/MC2/n108 ,
         \U1/aes_core/MC2/n107 , \U1/aes_core/MC2/n106 ,
         \U1/aes_core/MC2/n105 , \U1/aes_core/MC2/n104 ,
         \U1/aes_core/MC2/n103 , \U1/aes_core/MC2/n102 ,
         \U1/aes_core/MC2/n101 , \U1/aes_core/MC2/n100 , \U1/aes_core/MC2/n99 ,
         \U1/aes_core/MC2/n98 , \U1/aes_core/MC2/n97 , \U1/aes_core/MC2/n96 ,
         \U1/aes_core/MC2/n95 , \U1/aes_core/MC2/n94 , \U1/aes_core/MC2/n93 ,
         \U1/aes_core/MC2/n92 , \U1/aes_core/MC2/n91 , \U1/aes_core/MC2/n90 ,
         \U1/aes_core/MC2/n89 , \U1/aes_core/MC2/n88 , \U1/aes_core/MC2/n87 ,
         \U1/aes_core/MC2/n86 , \U1/aes_core/MC2/n85 , \U1/aes_core/MC2/n84 ,
         \U1/aes_core/MC2/n83 , \U1/aes_core/MC2/n82 , \U1/aes_core/MC2/n81 ,
         \U1/aes_core/MC2/n80 , \U1/aes_core/MC2/n79 , \U1/aes_core/MC2/n78 ,
         \U1/aes_core/MC2/n37 , \U1/aes_core/MC2/n34 , \U1/aes_core/MC2/n1 ,
         \U1/aes_core/MC3/n151 , \U1/aes_core/MC3/n150 ,
         \U1/aes_core/MC3/n149 , \U1/aes_core/MC3/n148 ,
         \U1/aes_core/MC3/n147 , \U1/aes_core/MC3/n146 ,
         \U1/aes_core/MC3/n145 , \U1/aes_core/MC3/n144 ,
         \U1/aes_core/MC3/n143 , \U1/aes_core/MC3/n142 ,
         \U1/aes_core/MC3/n141 , \U1/aes_core/MC3/n140 ,
         \U1/aes_core/MC3/n139 , \U1/aes_core/MC3/n138 ,
         \U1/aes_core/MC3/n137 , \U1/aes_core/MC3/n136 ,
         \U1/aes_core/MC3/n135 , \U1/aes_core/MC3/n134 ,
         \U1/aes_core/MC3/n133 , \U1/aes_core/MC3/n132 ,
         \U1/aes_core/MC3/n131 , \U1/aes_core/MC3/n130 ,
         \U1/aes_core/MC3/n129 , \U1/aes_core/MC3/n128 ,
         \U1/aes_core/MC3/n127 , \U1/aes_core/MC3/n126 ,
         \U1/aes_core/MC3/n125 , \U1/aes_core/MC3/n124 ,
         \U1/aes_core/MC3/n123 , \U1/aes_core/MC3/n122 ,
         \U1/aes_core/MC3/n121 , \U1/aes_core/MC3/n120 ,
         \U1/aes_core/MC3/n119 , \U1/aes_core/MC3/n118 ,
         \U1/aes_core/MC3/n117 , \U1/aes_core/MC3/n116 ,
         \U1/aes_core/MC3/n115 , \U1/aes_core/MC3/n114 ,
         \U1/aes_core/MC3/n113 , \U1/aes_core/MC3/n112 ,
         \U1/aes_core/MC3/n111 , \U1/aes_core/MC3/n110 ,
         \U1/aes_core/MC3/n109 , \U1/aes_core/MC3/n108 ,
         \U1/aes_core/MC3/n107 , \U1/aes_core/MC3/n106 ,
         \U1/aes_core/MC3/n105 , \U1/aes_core/MC3/n104 ,
         \U1/aes_core/MC3/n103 , \U1/aes_core/MC3/n102 ,
         \U1/aes_core/MC3/n101 , \U1/aes_core/MC3/n100 , \U1/aes_core/MC3/n99 ,
         \U1/aes_core/MC3/n98 , \U1/aes_core/MC3/n97 , \U1/aes_core/MC3/n96 ,
         \U1/aes_core/MC3/n95 , \U1/aes_core/MC3/n94 , \U1/aes_core/MC3/n93 ,
         \U1/aes_core/MC3/n92 , \U1/aes_core/MC3/n91 , \U1/aes_core/MC3/n90 ,
         \U1/aes_core/MC3/n89 , \U1/aes_core/MC3/n88 , \U1/aes_core/MC3/n87 ,
         \U1/aes_core/MC3/n86 , \U1/aes_core/MC3/n85 , \U1/aes_core/MC3/n84 ,
         \U1/aes_core/MC3/n83 , \U1/aes_core/MC3/n82 , \U1/aes_core/MC3/n81 ,
         \U1/aes_core/MC3/n80 , \U1/aes_core/MC3/n79 , \U1/aes_core/MC3/n78 ,
         \U1/aes_core/MC3/n37 , \U1/aes_core/MC3/n34 , \U1/aes_core/MC3/n1 ,
         \U1/keyexpantion/n8 , \U1/keyexpantion/n7 , \U1/keyexpantion/n6 ,
         \U1/keyexpantion/n5 , \U1/keyexpantion/n4 , \U1/keyexpantion/n3 ,
         \U1/keyexpantion/n2 , \U1/keyexpantion/n1 ,
         \U1/keyexpantion/SB0/n3362 , \U1/keyexpantion/SB0/n3361 ,
         \U1/keyexpantion/SB0/n3360 , \U1/keyexpantion/SB0/n3359 ,
         \U1/keyexpantion/SB0/n3358 , \U1/keyexpantion/SB0/n3357 ,
         \U1/keyexpantion/SB0/n3356 , \U1/keyexpantion/SB0/n3355 ,
         \U1/keyexpantion/SB0/n3354 , \U1/keyexpantion/SB0/n3353 ,
         \U1/keyexpantion/SB0/n3352 , \U1/keyexpantion/SB0/n3351 ,
         \U1/keyexpantion/SB0/n3350 , \U1/keyexpantion/SB0/n3349 ,
         \U1/keyexpantion/SB0/n3348 , \U1/keyexpantion/SB0/n3347 ,
         \U1/keyexpantion/SB0/n3346 , \U1/keyexpantion/SB0/n3345 ,
         \U1/keyexpantion/SB0/n3344 , \U1/keyexpantion/SB0/n3343 ,
         \U1/keyexpantion/SB0/n3342 , \U1/keyexpantion/SB0/n3341 ,
         \U1/keyexpantion/SB0/n3340 , \U1/keyexpantion/SB0/n3339 ,
         \U1/keyexpantion/SB0/n3338 , \U1/keyexpantion/SB0/n3337 ,
         \U1/keyexpantion/SB0/n3336 , \U1/keyexpantion/SB0/n3335 ,
         \U1/keyexpantion/SB0/n3334 , \U1/keyexpantion/SB0/n3333 ,
         \U1/keyexpantion/SB0/n3332 , \U1/keyexpantion/SB0/n3331 ,
         \U1/keyexpantion/SB0/n3330 , \U1/keyexpantion/SB0/n3329 ,
         \U1/keyexpantion/SB0/n3328 , \U1/keyexpantion/SB0/n3327 ,
         \U1/keyexpantion/SB0/n3326 , \U1/keyexpantion/SB0/n3325 ,
         \U1/keyexpantion/SB0/n3324 , \U1/keyexpantion/SB0/n3323 ,
         \U1/keyexpantion/SB0/n3322 , \U1/keyexpantion/SB0/n3321 ,
         \U1/keyexpantion/SB0/n3320 , \U1/keyexpantion/SB0/n3319 ,
         \U1/keyexpantion/SB0/n3318 , \U1/keyexpantion/SB0/n3317 ,
         \U1/keyexpantion/SB0/n3316 , \U1/keyexpantion/SB0/n3315 ,
         \U1/keyexpantion/SB0/n3314 , \U1/keyexpantion/SB0/n3313 ,
         \U1/keyexpantion/SB0/n3312 , \U1/keyexpantion/SB0/n3311 ,
         \U1/keyexpantion/SB0/n3310 , \U1/keyexpantion/SB0/n3309 ,
         \U1/keyexpantion/SB0/n3308 , \U1/keyexpantion/SB0/n3307 ,
         \U1/keyexpantion/SB0/n3306 , \U1/keyexpantion/SB0/n3305 ,
         \U1/keyexpantion/SB0/n3304 , \U1/keyexpantion/SB0/n3303 ,
         \U1/keyexpantion/SB0/n3302 , \U1/keyexpantion/SB0/n3301 ,
         \U1/keyexpantion/SB0/n3300 , \U1/keyexpantion/SB0/n3299 ,
         \U1/keyexpantion/SB0/n3298 , \U1/keyexpantion/SB0/n3297 ,
         \U1/keyexpantion/SB0/n3296 , \U1/keyexpantion/SB0/n3295 ,
         \U1/keyexpantion/SB0/n3294 , \U1/keyexpantion/SB0/n3293 ,
         \U1/keyexpantion/SB0/n3292 , \U1/keyexpantion/SB0/n3291 ,
         \U1/keyexpantion/SB0/n3290 , \U1/keyexpantion/SB0/n3289 ,
         \U1/keyexpantion/SB0/n3288 , \U1/keyexpantion/SB0/n3287 ,
         \U1/keyexpantion/SB0/n3286 , \U1/keyexpantion/SB0/n3285 ,
         \U1/keyexpantion/SB0/n3284 , \U1/keyexpantion/SB0/n3283 ,
         \U1/keyexpantion/SB0/n3282 , \U1/keyexpantion/SB0/n3281 ,
         \U1/keyexpantion/SB0/n3280 , \U1/keyexpantion/SB0/n3279 ,
         \U1/keyexpantion/SB0/n3278 , \U1/keyexpantion/SB0/n3277 ,
         \U1/keyexpantion/SB0/n3276 , \U1/keyexpantion/SB0/n3275 ,
         \U1/keyexpantion/SB0/n3274 , \U1/keyexpantion/SB0/n3273 ,
         \U1/keyexpantion/SB0/n3272 , \U1/keyexpantion/SB0/n3271 ,
         \U1/keyexpantion/SB0/n3270 , \U1/keyexpantion/SB0/n3269 ,
         \U1/keyexpantion/SB0/n3268 , \U1/keyexpantion/SB0/n3267 ,
         \U1/keyexpantion/SB0/n3266 , \U1/keyexpantion/SB0/n3265 ,
         \U1/keyexpantion/SB0/n3264 , \U1/keyexpantion/SB0/n3263 ,
         \U1/keyexpantion/SB0/n3262 , \U1/keyexpantion/SB0/n3261 ,
         \U1/keyexpantion/SB0/n3260 , \U1/keyexpantion/SB0/n3259 ,
         \U1/keyexpantion/SB0/n3258 , \U1/keyexpantion/SB0/n3257 ,
         \U1/keyexpantion/SB0/n3256 , \U1/keyexpantion/SB0/n3255 ,
         \U1/keyexpantion/SB0/n3254 , \U1/keyexpantion/SB0/n3253 ,
         \U1/keyexpantion/SB0/n3252 , \U1/keyexpantion/SB0/n3251 ,
         \U1/keyexpantion/SB0/n3250 , \U1/keyexpantion/SB0/n3249 ,
         \U1/keyexpantion/SB0/n3248 , \U1/keyexpantion/SB0/n3247 ,
         \U1/keyexpantion/SB0/n3246 , \U1/keyexpantion/SB0/n3245 ,
         \U1/keyexpantion/SB0/n3244 , \U1/keyexpantion/SB0/n3243 ,
         \U1/keyexpantion/SB0/n3242 , \U1/keyexpantion/SB0/n3241 ,
         \U1/keyexpantion/SB0/n3240 , \U1/keyexpantion/SB0/n3239 ,
         \U1/keyexpantion/SB0/n3238 , \U1/keyexpantion/SB0/n3237 ,
         \U1/keyexpantion/SB0/n3236 , \U1/keyexpantion/SB0/n3235 ,
         \U1/keyexpantion/SB0/n3234 , \U1/keyexpantion/SB0/n3233 ,
         \U1/keyexpantion/SB0/n3232 , \U1/keyexpantion/SB0/n3231 ,
         \U1/keyexpantion/SB0/n3230 , \U1/keyexpantion/SB0/n3229 ,
         \U1/keyexpantion/SB0/n3228 , \U1/keyexpantion/SB0/n3227 ,
         \U1/keyexpantion/SB0/n3226 , \U1/keyexpantion/SB0/n3225 ,
         \U1/keyexpantion/SB0/n3224 , \U1/keyexpantion/SB0/n3223 ,
         \U1/keyexpantion/SB0/n3222 , \U1/keyexpantion/SB0/n3221 ,
         \U1/keyexpantion/SB0/n3220 , \U1/keyexpantion/SB0/n3219 ,
         \U1/keyexpantion/SB0/n3218 , \U1/keyexpantion/SB0/n3217 ,
         \U1/keyexpantion/SB0/n3216 , \U1/keyexpantion/SB0/n3215 ,
         \U1/keyexpantion/SB0/n3214 , \U1/keyexpantion/SB0/n3213 ,
         \U1/keyexpantion/SB0/n3212 , \U1/keyexpantion/SB0/n3211 ,
         \U1/keyexpantion/SB0/n3210 , \U1/keyexpantion/SB0/n3209 ,
         \U1/keyexpantion/SB0/n3208 , \U1/keyexpantion/SB0/n3207 ,
         \U1/keyexpantion/SB0/n3206 , \U1/keyexpantion/SB0/n3205 ,
         \U1/keyexpantion/SB0/n3204 , \U1/keyexpantion/SB0/n3203 ,
         \U1/keyexpantion/SB0/n3202 , \U1/keyexpantion/SB0/n3201 ,
         \U1/keyexpantion/SB0/n3200 , \U1/keyexpantion/SB0/n3199 ,
         \U1/keyexpantion/SB0/n3198 , \U1/keyexpantion/SB0/n3197 ,
         \U1/keyexpantion/SB0/n3196 , \U1/keyexpantion/SB0/n3195 ,
         \U1/keyexpantion/SB0/n3194 , \U1/keyexpantion/SB0/n3193 ,
         \U1/keyexpantion/SB0/n3192 , \U1/keyexpantion/SB0/n3191 ,
         \U1/keyexpantion/SB0/n3190 , \U1/keyexpantion/SB0/n3189 ,
         \U1/keyexpantion/SB0/n3188 , \U1/keyexpantion/SB0/n3187 ,
         \U1/keyexpantion/SB0/n3186 , \U1/keyexpantion/SB0/n3185 ,
         \U1/keyexpantion/SB0/n3184 , \U1/keyexpantion/SB0/n3183 ,
         \U1/keyexpantion/SB0/n3182 , \U1/keyexpantion/SB0/n3181 ,
         \U1/keyexpantion/SB0/n3180 , \U1/keyexpantion/SB0/n3179 ,
         \U1/keyexpantion/SB0/n3178 , \U1/keyexpantion/SB0/n3177 ,
         \U1/keyexpantion/SB0/n3176 , \U1/keyexpantion/SB0/n3175 ,
         \U1/keyexpantion/SB0/n3174 , \U1/keyexpantion/SB0/n3173 ,
         \U1/keyexpantion/SB0/n3172 , \U1/keyexpantion/SB0/n3171 ,
         \U1/keyexpantion/SB0/n3170 , \U1/keyexpantion/SB0/n3169 ,
         \U1/keyexpantion/SB0/n3168 , \U1/keyexpantion/SB0/n3167 ,
         \U1/keyexpantion/SB0/n3166 , \U1/keyexpantion/SB0/n3165 ,
         \U1/keyexpantion/SB0/n3164 , \U1/keyexpantion/SB0/n3163 ,
         \U1/keyexpantion/SB0/n3162 , \U1/keyexpantion/SB0/n3161 ,
         \U1/keyexpantion/SB0/n3160 , \U1/keyexpantion/SB0/n3159 ,
         \U1/keyexpantion/SB0/n3158 , \U1/keyexpantion/SB0/n3157 ,
         \U1/keyexpantion/SB0/n3156 , \U1/keyexpantion/SB0/n3155 ,
         \U1/keyexpantion/SB0/n3154 , \U1/keyexpantion/SB0/n3153 ,
         \U1/keyexpantion/SB0/n3152 , \U1/keyexpantion/SB0/n3151 ,
         \U1/keyexpantion/SB0/n3150 , \U1/keyexpantion/SB0/n3149 ,
         \U1/keyexpantion/SB0/n3148 , \U1/keyexpantion/SB0/n3147 ,
         \U1/keyexpantion/SB0/n3146 , \U1/keyexpantion/SB0/n3145 ,
         \U1/keyexpantion/SB0/n3144 , \U1/keyexpantion/SB0/n3143 ,
         \U1/keyexpantion/SB0/n3142 , \U1/keyexpantion/SB0/n3141 ,
         \U1/keyexpantion/SB0/n3140 , \U1/keyexpantion/SB0/n3139 ,
         \U1/keyexpantion/SB0/n3138 , \U1/keyexpantion/SB0/n3137 ,
         \U1/keyexpantion/SB0/n3136 , \U1/keyexpantion/SB0/n3135 ,
         \U1/keyexpantion/SB0/n3134 , \U1/keyexpantion/SB0/n3133 ,
         \U1/keyexpantion/SB0/n3132 , \U1/keyexpantion/SB0/n3131 ,
         \U1/keyexpantion/SB0/n3130 , \U1/keyexpantion/SB0/n3129 ,
         \U1/keyexpantion/SB0/n3128 , \U1/keyexpantion/SB0/n3127 ,
         \U1/keyexpantion/SB0/n3126 , \U1/keyexpantion/SB0/n3125 ,
         \U1/keyexpantion/SB0/n3124 , \U1/keyexpantion/SB0/n3123 ,
         \U1/keyexpantion/SB0/n3122 , \U1/keyexpantion/SB0/n3121 ,
         \U1/keyexpantion/SB0/n3120 , \U1/keyexpantion/SB0/n3119 ,
         \U1/keyexpantion/SB0/n3118 , \U1/keyexpantion/SB0/n3117 ,
         \U1/keyexpantion/SB0/n3116 , \U1/keyexpantion/SB0/n3115 ,
         \U1/keyexpantion/SB0/n3114 , \U1/keyexpantion/SB0/n3113 ,
         \U1/keyexpantion/SB0/n3112 , \U1/keyexpantion/SB0/n3111 ,
         \U1/keyexpantion/SB0/n3110 , \U1/keyexpantion/SB0/n3109 ,
         \U1/keyexpantion/SB0/n3108 , \U1/keyexpantion/SB0/n3107 ,
         \U1/keyexpantion/SB0/n3106 , \U1/keyexpantion/SB0/n3105 ,
         \U1/keyexpantion/SB0/n3104 , \U1/keyexpantion/SB0/n3103 ,
         \U1/keyexpantion/SB0/n3102 , \U1/keyexpantion/SB0/n3101 ,
         \U1/keyexpantion/SB0/n3100 , \U1/keyexpantion/SB0/n3099 ,
         \U1/keyexpantion/SB0/n3098 , \U1/keyexpantion/SB0/n3097 ,
         \U1/keyexpantion/SB0/n3096 , \U1/keyexpantion/SB0/n3095 ,
         \U1/keyexpantion/SB0/n3094 , \U1/keyexpantion/SB0/n3093 ,
         \U1/keyexpantion/SB0/n3092 , \U1/keyexpantion/SB0/n3091 ,
         \U1/keyexpantion/SB0/n3090 , \U1/keyexpantion/SB0/n3089 ,
         \U1/keyexpantion/SB0/n3088 , \U1/keyexpantion/SB0/n3087 ,
         \U1/keyexpantion/SB0/n3086 , \U1/keyexpantion/SB0/n3085 ,
         \U1/keyexpantion/SB0/n3084 , \U1/keyexpantion/SB0/n3083 ,
         \U1/keyexpantion/SB0/n3082 , \U1/keyexpantion/SB0/n3081 ,
         \U1/keyexpantion/SB0/n3080 , \U1/keyexpantion/SB0/n3079 ,
         \U1/keyexpantion/SB0/n3078 , \U1/keyexpantion/SB0/n3077 ,
         \U1/keyexpantion/SB0/n3076 , \U1/keyexpantion/SB0/n3075 ,
         \U1/keyexpantion/SB0/n3074 , \U1/keyexpantion/SB0/n3073 ,
         \U1/keyexpantion/SB0/n3072 , \U1/keyexpantion/SB0/n3071 ,
         \U1/keyexpantion/SB0/n3070 , \U1/keyexpantion/SB0/n3069 ,
         \U1/keyexpantion/SB0/n3068 , \U1/keyexpantion/SB0/n3067 ,
         \U1/keyexpantion/SB0/n3066 , \U1/keyexpantion/SB0/n3065 ,
         \U1/keyexpantion/SB0/n3064 , \U1/keyexpantion/SB0/n3063 ,
         \U1/keyexpantion/SB0/n3062 , \U1/keyexpantion/SB0/n3061 ,
         \U1/keyexpantion/SB0/n3060 , \U1/keyexpantion/SB0/n3059 ,
         \U1/keyexpantion/SB0/n3058 , \U1/keyexpantion/SB0/n3057 ,
         \U1/keyexpantion/SB0/n3056 , \U1/keyexpantion/SB0/n3055 ,
         \U1/keyexpantion/SB0/n3054 , \U1/keyexpantion/SB0/n3053 ,
         \U1/keyexpantion/SB0/n3052 , \U1/keyexpantion/SB0/n3051 ,
         \U1/keyexpantion/SB0/n3050 , \U1/keyexpantion/SB0/n3049 ,
         \U1/keyexpantion/SB0/n3048 , \U1/keyexpantion/SB0/n3047 ,
         \U1/keyexpantion/SB0/n3046 , \U1/keyexpantion/SB0/n3045 ,
         \U1/keyexpantion/SB0/n3044 , \U1/keyexpantion/SB0/n3043 ,
         \U1/keyexpantion/SB0/n3042 , \U1/keyexpantion/SB0/n3041 ,
         \U1/keyexpantion/SB0/n3040 , \U1/keyexpantion/SB0/n3039 ,
         \U1/keyexpantion/SB0/n3038 , \U1/keyexpantion/SB0/n3037 ,
         \U1/keyexpantion/SB0/n3036 , \U1/keyexpantion/SB0/n3035 ,
         \U1/keyexpantion/SB0/n3034 , \U1/keyexpantion/SB0/n3033 ,
         \U1/keyexpantion/SB0/n3032 , \U1/keyexpantion/SB0/n3031 ,
         \U1/keyexpantion/SB0/n3030 , \U1/keyexpantion/SB0/n3029 ,
         \U1/keyexpantion/SB0/n3028 , \U1/keyexpantion/SB0/n3027 ,
         \U1/keyexpantion/SB0/n3026 , \U1/keyexpantion/SB0/n3025 ,
         \U1/keyexpantion/SB0/n3024 , \U1/keyexpantion/SB0/n3023 ,
         \U1/keyexpantion/SB0/n3022 , \U1/keyexpantion/SB0/n3021 ,
         \U1/keyexpantion/SB0/n3020 , \U1/keyexpantion/SB0/n3019 ,
         \U1/keyexpantion/SB0/n3018 , \U1/keyexpantion/SB0/n3017 ,
         \U1/keyexpantion/SB0/n3016 , \U1/keyexpantion/SB0/n3015 ,
         \U1/keyexpantion/SB0/n3014 , \U1/keyexpantion/SB0/n3013 ,
         \U1/keyexpantion/SB0/n3012 , \U1/keyexpantion/SB0/n3011 ,
         \U1/keyexpantion/SB0/n3010 , \U1/keyexpantion/SB0/n3009 ,
         \U1/keyexpantion/SB0/n3008 , \U1/keyexpantion/SB0/n3007 ,
         \U1/keyexpantion/SB0/n3006 , \U1/keyexpantion/SB0/n3005 ,
         \U1/keyexpantion/SB0/n3004 , \U1/keyexpantion/SB0/n3003 ,
         \U1/keyexpantion/SB0/n3002 , \U1/keyexpantion/SB0/n3001 ,
         \U1/keyexpantion/SB0/n3000 , \U1/keyexpantion/SB0/n2999 ,
         \U1/keyexpantion/SB0/n2998 , \U1/keyexpantion/SB0/n2997 ,
         \U1/keyexpantion/SB0/n2996 , \U1/keyexpantion/SB0/n2995 ,
         \U1/keyexpantion/SB0/n2994 , \U1/keyexpantion/SB0/n2993 ,
         \U1/keyexpantion/SB0/n2992 , \U1/keyexpantion/SB0/n2991 ,
         \U1/keyexpantion/SB0/n2990 , \U1/keyexpantion/SB0/n2989 ,
         \U1/keyexpantion/SB0/n2988 , \U1/keyexpantion/SB0/n2987 ,
         \U1/keyexpantion/SB0/n2986 , \U1/keyexpantion/SB0/n2985 ,
         \U1/keyexpantion/SB0/n2984 , \U1/keyexpantion/SB0/n2983 ,
         \U1/keyexpantion/SB0/n2982 , \U1/keyexpantion/SB0/n2981 ,
         \U1/keyexpantion/SB0/n2980 , \U1/keyexpantion/SB0/n2979 ,
         \U1/keyexpantion/SB0/n2978 , \U1/keyexpantion/SB0/n2977 ,
         \U1/keyexpantion/SB0/n2976 , \U1/keyexpantion/SB0/n2975 ,
         \U1/keyexpantion/SB0/n2974 , \U1/keyexpantion/SB0/n2973 ,
         \U1/keyexpantion/SB0/n2972 , \U1/keyexpantion/SB0/n2971 ,
         \U1/keyexpantion/SB0/n2970 , \U1/keyexpantion/SB0/n2969 ,
         \U1/keyexpantion/SB0/n2968 , \U1/keyexpantion/SB0/n2967 ,
         \U1/keyexpantion/SB0/n2966 , \U1/keyexpantion/SB0/n2965 ,
         \U1/keyexpantion/SB0/n2964 , \U1/keyexpantion/SB0/n2963 ,
         \U1/keyexpantion/SB0/n2962 , \U1/keyexpantion/SB0/n2961 ,
         \U1/keyexpantion/SB0/n2960 , \U1/keyexpantion/SB0/n2959 ,
         \U1/keyexpantion/SB0/n2958 , \U1/keyexpantion/SB0/n2957 ,
         \U1/keyexpantion/SB0/n2956 , \U1/keyexpantion/SB0/n2955 ,
         \U1/keyexpantion/SB0/n2954 , \U1/keyexpantion/SB0/n2953 ,
         \U1/keyexpantion/SB0/n2952 , \U1/keyexpantion/SB0/n2951 ,
         \U1/keyexpantion/SB0/n2950 , \U1/keyexpantion/SB0/n2949 ,
         \U1/keyexpantion/SB0/n2948 , \U1/keyexpantion/SB0/n2947 ,
         \U1/keyexpantion/SB0/n2946 , \U1/keyexpantion/SB0/n2945 ,
         \U1/keyexpantion/SB0/n2944 , \U1/keyexpantion/SB0/n2943 ,
         \U1/keyexpantion/SB0/n2942 , \U1/keyexpantion/SB0/n2941 ,
         \U1/keyexpantion/SB0/n2940 , \U1/keyexpantion/SB0/n2939 ,
         \U1/keyexpantion/SB0/n2938 , \U1/keyexpantion/SB0/n2937 ,
         \U1/keyexpantion/SB0/n2936 , \U1/keyexpantion/SB0/n2935 ,
         \U1/keyexpantion/SB0/n2934 , \U1/keyexpantion/SB0/n2933 ,
         \U1/keyexpantion/SB0/n2932 , \U1/keyexpantion/SB0/n2931 ,
         \U1/keyexpantion/SB0/n2930 , \U1/keyexpantion/SB0/n2929 ,
         \U1/keyexpantion/SB0/n2928 , \U1/keyexpantion/SB0/n2927 ,
         \U1/keyexpantion/SB0/n2926 , \U1/keyexpantion/SB0/n2925 ,
         \U1/keyexpantion/SB0/n2924 , \U1/keyexpantion/SB0/n2923 ,
         \U1/keyexpantion/SB0/n2922 , \U1/keyexpantion/SB0/n2921 ,
         \U1/keyexpantion/SB0/n2920 , \U1/keyexpantion/SB0/n2919 ,
         \U1/keyexpantion/SB0/n2918 , \U1/keyexpantion/SB0/n2917 ,
         \U1/keyexpantion/SB0/n2916 , \U1/keyexpantion/SB0/n2915 ,
         \U1/keyexpantion/SB0/n2914 , \U1/keyexpantion/SB0/n2913 ,
         \U1/keyexpantion/SB0/n2912 , \U1/keyexpantion/SB0/n2911 ,
         \U1/keyexpantion/SB0/n2910 , \U1/keyexpantion/SB0/n2909 ,
         \U1/keyexpantion/SB0/n2908 , \U1/keyexpantion/SB0/n2907 ,
         \U1/keyexpantion/SB0/n2906 , \U1/keyexpantion/SB0/n2905 ,
         \U1/keyexpantion/SB0/n2904 , \U1/keyexpantion/SB0/n2903 ,
         \U1/keyexpantion/SB0/n2902 , \U1/keyexpantion/SB0/n2901 ,
         \U1/keyexpantion/SB0/n2900 , \U1/keyexpantion/SB0/n2899 ,
         \U1/keyexpantion/SB0/n2898 , \U1/keyexpantion/SB0/n2897 ,
         \U1/keyexpantion/SB0/n2896 , \U1/keyexpantion/SB0/n2895 ,
         \U1/keyexpantion/SB0/n2894 , \U1/keyexpantion/SB0/n2893 ,
         \U1/keyexpantion/SB0/n2892 , \U1/keyexpantion/SB0/n2891 ,
         \U1/keyexpantion/SB0/n2890 , \U1/keyexpantion/SB0/n2889 ,
         \U1/keyexpantion/SB0/n2888 , \U1/keyexpantion/SB0/n2887 ,
         \U1/keyexpantion/SB0/n2886 , \U1/keyexpantion/SB0/n2885 ,
         \U1/keyexpantion/SB0/n2884 , \U1/keyexpantion/SB0/n2883 ,
         \U1/keyexpantion/SB0/n2882 , \U1/keyexpantion/SB0/n2881 ,
         \U1/keyexpantion/SB0/n2880 , \U1/keyexpantion/SB0/n2879 ,
         \U1/keyexpantion/SB0/n2878 , \U1/keyexpantion/SB0/n2877 ,
         \U1/keyexpantion/SB0/n2876 , \U1/keyexpantion/SB0/n2875 ,
         \U1/keyexpantion/SB0/n2874 , \U1/keyexpantion/SB0/n2873 ,
         \U1/keyexpantion/SB0/n2872 , \U1/keyexpantion/SB0/n2871 ,
         \U1/keyexpantion/SB0/n2870 , \U1/keyexpantion/SB0/n2869 ,
         \U1/keyexpantion/SB0/n2868 , \U1/keyexpantion/SB0/n2867 ,
         \U1/keyexpantion/SB0/n2866 , \U1/keyexpantion/SB0/n2865 ,
         \U1/keyexpantion/SB0/n2864 , \U1/keyexpantion/SB0/n2863 ,
         \U1/keyexpantion/SB0/n2862 , \U1/keyexpantion/SB0/n2861 ,
         \U1/keyexpantion/SB0/n2860 , \U1/keyexpantion/SB0/n2859 ,
         \U1/keyexpantion/SB0/n2858 , \U1/keyexpantion/SB0/n2857 ,
         \U1/keyexpantion/SB0/n2856 , \U1/keyexpantion/SB0/n2855 ,
         \U1/keyexpantion/SB0/n2854 , \U1/keyexpantion/SB0/n2853 ,
         \U1/keyexpantion/SB0/n2852 , \U1/keyexpantion/SB0/n2851 ,
         \U1/keyexpantion/SB0/n2850 , \U1/keyexpantion/SB0/n2849 ,
         \U1/keyexpantion/SB0/n2848 , \U1/keyexpantion/SB0/n2847 ,
         \U1/keyexpantion/SB0/n2846 , \U1/keyexpantion/SB0/n2845 ,
         \U1/keyexpantion/SB0/n2844 , \U1/keyexpantion/SB0/n2843 ,
         \U1/keyexpantion/SB0/n2842 , \U1/keyexpantion/SB0/n2841 ,
         \U1/keyexpantion/SB0/n2840 , \U1/keyexpantion/SB0/n2839 ,
         \U1/keyexpantion/SB0/n2838 , \U1/keyexpantion/SB0/n2837 ,
         \U1/keyexpantion/SB0/n2836 , \U1/keyexpantion/SB0/n2835 ,
         \U1/keyexpantion/SB0/n2834 , \U1/keyexpantion/SB0/n2833 ,
         \U1/keyexpantion/SB0/n2832 , \U1/keyexpantion/SB0/n2831 ,
         \U1/keyexpantion/SB0/n2830 , \U1/keyexpantion/SB0/n2829 ,
         \U1/keyexpantion/SB0/n2828 , \U1/keyexpantion/SB0/n2827 ,
         \U1/keyexpantion/SB0/n2826 , \U1/keyexpantion/SB0/n2825 ,
         \U1/keyexpantion/SB0/n2824 , \U1/keyexpantion/SB0/n2823 ,
         \U1/keyexpantion/SB0/n2822 , \U1/keyexpantion/SB0/n2821 ,
         \U1/keyexpantion/SB0/n2820 , \U1/keyexpantion/SB0/n2819 ,
         \U1/keyexpantion/SB0/n2818 , \U1/keyexpantion/SB0/n2817 ,
         \U1/keyexpantion/SB0/n2816 , \U1/keyexpantion/SB0/n2815 ,
         \U1/keyexpantion/SB0/n2814 , \U1/keyexpantion/SB0/n2813 ,
         \U1/keyexpantion/SB0/n2812 , \U1/keyexpantion/SB0/n2811 ,
         \U1/keyexpantion/SB0/n2810 , \U1/keyexpantion/SB0/n2809 ,
         \U1/keyexpantion/SB0/n2808 , \U1/keyexpantion/SB0/n2807 ,
         \U1/keyexpantion/SB0/n2806 , \U1/keyexpantion/SB0/n2805 ,
         \U1/keyexpantion/SB0/n2804 , \U1/keyexpantion/SB0/n2803 ,
         \U1/keyexpantion/SB0/n2802 , \U1/keyexpantion/SB0/n2801 ,
         \U1/keyexpantion/SB0/n2800 , \U1/keyexpantion/SB0/n2799 ,
         \U1/keyexpantion/SB0/n2798 , \U1/keyexpantion/SB0/n2797 ,
         \U1/keyexpantion/SB0/n2796 , \U1/keyexpantion/SB0/n2795 ,
         \U1/keyexpantion/SB0/n2794 , \U1/keyexpantion/SB0/n2793 ,
         \U1/keyexpantion/SB0/n2792 , \U1/keyexpantion/SB0/n2791 ,
         \U1/keyexpantion/SB0/n2790 , \U1/keyexpantion/SB0/n2789 ,
         \U1/keyexpantion/SB0/n2788 , \U1/keyexpantion/SB0/n2787 ,
         \U1/keyexpantion/SB0/n2786 , \U1/keyexpantion/SB0/n2785 ,
         \U1/keyexpantion/SB0/n2784 , \U1/keyexpantion/SB0/n2783 ,
         \U1/keyexpantion/SB0/n2782 , \U1/keyexpantion/SB0/n2781 ,
         \U1/keyexpantion/SB0/n2780 , \U1/keyexpantion/SB0/n2779 ,
         \U1/keyexpantion/SB0/n2778 , \U1/keyexpantion/SB0/n2777 ,
         \U1/keyexpantion/SB0/n2776 , \U1/keyexpantion/SB0/n2775 ,
         \U1/keyexpantion/SB0/n2774 , \U1/keyexpantion/SB0/n2773 ,
         \U1/keyexpantion/SB0/n2772 , \U1/keyexpantion/SB0/n2771 ,
         \U1/keyexpantion/SB0/n2770 , \U1/keyexpantion/SB0/n2769 ,
         \U1/keyexpantion/SB0/n2768 , \U1/keyexpantion/SB0/n2767 ,
         \U1/keyexpantion/SB0/n2766 , \U1/keyexpantion/SB0/n2765 ,
         \U1/keyexpantion/SB0/n2764 , \U1/keyexpantion/SB0/n2763 ,
         \U1/keyexpantion/SB0/n2762 , \U1/keyexpantion/SB0/n2761 ,
         \U1/keyexpantion/SB0/n2760 , \U1/keyexpantion/SB0/n2759 ,
         \U1/keyexpantion/SB0/n2758 , \U1/keyexpantion/SB0/n2757 ,
         \U1/keyexpantion/SB0/n2756 , \U1/keyexpantion/SB0/n2755 ,
         \U1/keyexpantion/SB0/n2754 , \U1/keyexpantion/SB0/n2753 ,
         \U1/keyexpantion/SB0/n2752 , \U1/keyexpantion/SB0/n2751 ,
         \U1/keyexpantion/SB0/n2750 , \U1/keyexpantion/SB0/n2749 ,
         \U1/keyexpantion/SB0/n2748 , \U1/keyexpantion/SB0/n2747 ,
         \U1/keyexpantion/SB0/n2746 , \U1/keyexpantion/SB0/n2745 ,
         \U1/keyexpantion/SB0/n2744 , \U1/keyexpantion/SB0/n2743 ,
         \U1/keyexpantion/SB0/n2742 , \U1/keyexpantion/SB0/n2741 ,
         \U1/keyexpantion/SB0/n2740 , \U1/keyexpantion/SB0/n2739 ,
         \U1/keyexpantion/SB0/n2738 , \U1/keyexpantion/SB0/n2737 ,
         \U1/keyexpantion/SB0/n2736 , \U1/keyexpantion/SB0/n2735 ,
         \U1/keyexpantion/SB0/n2734 , \U1/keyexpantion/SB0/n2733 ,
         \U1/keyexpantion/SB0/n2732 , \U1/keyexpantion/SB0/n2731 ,
         \U1/keyexpantion/SB0/n2730 , \U1/keyexpantion/SB0/n2729 ,
         \U1/keyexpantion/SB0/n2728 , \U1/keyexpantion/SB0/n2727 ,
         \U1/keyexpantion/SB0/n2726 , \U1/keyexpantion/SB0/n2725 ,
         \U1/keyexpantion/SB0/n2724 , \U1/keyexpantion/SB0/n2723 ,
         \U1/keyexpantion/SB0/n2722 , \U1/keyexpantion/SB0/n2721 ,
         \U1/keyexpantion/SB0/n2720 , \U1/keyexpantion/SB0/n2719 ,
         \U1/keyexpantion/SB0/n2718 , \U1/keyexpantion/SB0/n2717 ,
         \U1/keyexpantion/SB0/n2716 , \U1/keyexpantion/SB0/n2715 ,
         \U1/keyexpantion/SB0/n2714 , \U1/keyexpantion/SB0/n2713 ,
         \U1/keyexpantion/SB0/n2712 , \U1/keyexpantion/SB0/n2711 ,
         \U1/keyexpantion/SB0/n2710 , \U1/keyexpantion/SB0/n2709 ,
         \U1/keyexpantion/SB0/n2708 , \U1/keyexpantion/SB0/n2707 ,
         \U1/keyexpantion/SB0/n2706 , \U1/keyexpantion/SB0/n2705 ,
         \U1/keyexpantion/SB0/n2704 , \U1/keyexpantion/SB0/n2703 ,
         \U1/keyexpantion/SB0/n2702 , \U1/keyexpantion/SB0/n2701 ,
         \U1/keyexpantion/SB0/n2700 , \U1/keyexpantion/SB0/n2699 ,
         \U1/keyexpantion/SB0/n2698 , \U1/keyexpantion/SB0/n2697 ,
         \U1/keyexpantion/SB0/n2696 , \U1/keyexpantion/SB0/n2695 ,
         \U1/keyexpantion/SB0/n2694 , \U1/keyexpantion/SB0/n2693 ,
         \U1/keyexpantion/SB0/n2692 , \U1/keyexpantion/SB0/n2691 ,
         \U1/keyexpantion/SB0/n2690 , \U1/keyexpantion/SB0/n2689 ,
         \U1/keyexpantion/SB0/n2688 , \U1/keyexpantion/SB0/n2687 ,
         \U1/keyexpantion/SB0/n2686 , \U1/keyexpantion/SB0/n2685 ,
         \U1/keyexpantion/SB0/n2684 , \U1/keyexpantion/SB0/n2683 ,
         \U1/keyexpantion/SB0/n2682 , \U1/keyexpantion/SB0/n2681 ,
         \U1/keyexpantion/SB0/n2680 , \U1/keyexpantion/SB0/n2679 ,
         \U1/keyexpantion/SB0/n2678 , \U1/keyexpantion/SB0/n2677 ,
         \U1/keyexpantion/SB0/n2676 , \U1/keyexpantion/SB0/n2675 ,
         \U1/keyexpantion/SB0/n2674 , \U1/keyexpantion/SB0/n2673 ,
         \U1/keyexpantion/SB0/n2672 , \U1/keyexpantion/SB0/n2671 ,
         \U1/keyexpantion/SB0/n2670 , \U1/keyexpantion/SB0/n2669 ,
         \U1/keyexpantion/SB0/n2668 , \U1/keyexpantion/SB0/n2667 ,
         \U1/keyexpantion/SB0/n2666 , \U1/keyexpantion/SB0/n2665 ,
         \U1/keyexpantion/SB0/n2664 , \U1/keyexpantion/SB0/n2663 ,
         \U1/keyexpantion/SB0/n2662 , \U1/keyexpantion/SB0/n2661 ,
         \U1/keyexpantion/SB0/n2660 , \U1/keyexpantion/SB0/n2659 ,
         \U1/keyexpantion/SB0/n2658 , \U1/keyexpantion/SB0/n2657 ,
         \U1/keyexpantion/SB0/n2656 , \U1/keyexpantion/SB0/n2655 ,
         \U1/keyexpantion/SB0/n2654 , \U1/keyexpantion/SB0/n2653 ,
         \U1/keyexpantion/SB0/n2652 , \U1/keyexpantion/SB0/n2651 ,
         \U1/keyexpantion/SB0/n2650 , \U1/keyexpantion/SB0/n2649 ,
         \U1/keyexpantion/SB0/n2648 , \U1/keyexpantion/SB0/n2647 ,
         \U1/keyexpantion/SB0/n2646 , \U1/keyexpantion/SB0/n2645 ,
         \U1/keyexpantion/SB0/n2644 , \U1/keyexpantion/SB0/n2643 ,
         \U1/keyexpantion/SB0/n2642 , \U1/keyexpantion/SB0/n2641 ,
         \U1/keyexpantion/SB0/n2640 , \U1/keyexpantion/SB0/n2639 ,
         \U1/keyexpantion/SB0/n2638 , \U1/keyexpantion/SB0/n2637 ,
         \U1/keyexpantion/SB0/n2636 , \U1/keyexpantion/SB0/n2635 ,
         \U1/keyexpantion/SB0/n2634 , \U1/keyexpantion/SB0/n2633 ,
         \U1/keyexpantion/SB0/n2632 , \U1/keyexpantion/SB0/n2631 ,
         \U1/keyexpantion/SB0/n2630 , \U1/keyexpantion/SB0/n2629 ,
         \U1/keyexpantion/SB0/n2628 , \U1/keyexpantion/SB0/n2627 ,
         \U1/keyexpantion/SB0/n2626 , \U1/keyexpantion/SB0/n2625 ,
         \U1/keyexpantion/SB0/n2624 , \U1/keyexpantion/SB0/n2623 ,
         \U1/keyexpantion/SB0/n2622 , \U1/keyexpantion/SB0/n2621 ,
         \U1/keyexpantion/SB0/n2620 , \U1/keyexpantion/SB0/n2619 ,
         \U1/keyexpantion/SB0/n2618 , \U1/keyexpantion/SB0/n2617 ,
         \U1/keyexpantion/SB0/n2616 , \U1/keyexpantion/SB0/n2615 ,
         \U1/keyexpantion/SB0/n2614 , \U1/keyexpantion/SB0/n2613 ,
         \U1/keyexpantion/SB0/n2612 , \U1/keyexpantion/SB0/n2611 ,
         \U1/keyexpantion/SB0/n2610 , \U1/keyexpantion/SB0/n2609 ,
         \U1/keyexpantion/SB0/n2608 , \U1/keyexpantion/SB0/n2607 ,
         \U1/keyexpantion/SB0/n2606 , \U1/keyexpantion/SB0/n2605 ,
         \U1/keyexpantion/SB0/n2604 , \U1/keyexpantion/SB0/n2603 ,
         \U1/keyexpantion/SB0/n2602 , \U1/keyexpantion/SB0/n2601 ,
         \U1/keyexpantion/SB0/n2600 , \U1/keyexpantion/SB0/n2599 ,
         \U1/keyexpantion/SB0/n2598 , \U1/keyexpantion/SB0/n2597 ,
         \U1/keyexpantion/SB0/n2596 , \U1/keyexpantion/SB0/n2595 ,
         \U1/keyexpantion/SB0/n2594 , \U1/keyexpantion/SB0/n2593 ,
         \U1/keyexpantion/SB0/n2592 , \U1/keyexpantion/SB0/n2591 ,
         \U1/keyexpantion/SB0/n2590 , \U1/keyexpantion/SB0/n2589 ,
         \U1/keyexpantion/SB0/n2588 , \U1/keyexpantion/SB0/n2587 ,
         \U1/keyexpantion/SB0/n2586 , \U1/keyexpantion/SB0/n2585 ,
         \U1/keyexpantion/SB0/n2584 , \U1/keyexpantion/SB0/n2583 ,
         \U1/keyexpantion/SB0/n2582 , \U1/keyexpantion/SB0/n2581 ,
         \U1/keyexpantion/SB0/n2580 , \U1/keyexpantion/SB0/n2579 ,
         \U1/keyexpantion/SB0/n2578 , \U1/keyexpantion/SB0/n2577 ,
         \U1/keyexpantion/SB0/n2576 , \U1/keyexpantion/SB0/n2575 ,
         \U1/keyexpantion/SB0/n2574 , \U1/keyexpantion/SB0/n2573 ,
         \U1/keyexpantion/SB0/n2572 , \U1/keyexpantion/SB0/n2571 ,
         \U1/keyexpantion/SB0/n2570 , \U1/keyexpantion/SB0/n2569 ,
         \U1/keyexpantion/SB0/n2568 , \U1/keyexpantion/SB0/n2567 ,
         \U1/keyexpantion/SB0/n2566 , \U1/keyexpantion/SB0/n2565 ,
         \U1/keyexpantion/SB0/n2564 , \U1/keyexpantion/SB0/n2563 ,
         \U1/keyexpantion/SB0/n2562 , \U1/keyexpantion/SB0/n2561 ,
         \U1/keyexpantion/SB0/n2560 , \U1/keyexpantion/SB0/n2559 ,
         \U1/keyexpantion/SB0/n2558 , \U1/keyexpantion/SB0/n2557 ,
         \U1/keyexpantion/SB0/n2556 , \U1/keyexpantion/SB0/n2555 ,
         \U1/keyexpantion/SB0/n2554 , \U1/keyexpantion/SB0/n2553 ,
         \U1/keyexpantion/SB0/n2552 , \U1/keyexpantion/SB0/n2551 ,
         \U1/keyexpantion/SB0/n2550 , \U1/keyexpantion/SB0/n2549 ,
         \U1/keyexpantion/SB0/n2548 , \U1/keyexpantion/SB0/n2547 ,
         \U1/keyexpantion/SB0/n2546 , \U1/keyexpantion/SB0/n2545 ,
         \U1/keyexpantion/SB0/n2544 , \U1/keyexpantion/SB0/n2543 ,
         \U1/keyexpantion/SB0/n2542 , \U1/keyexpantion/SB0/n2541 ,
         \U1/keyexpantion/SB0/n2540 , \U1/keyexpantion/SB0/n2539 ,
         \U1/keyexpantion/SB0/n2538 , \U1/keyexpantion/SB0/n2537 ,
         \U1/keyexpantion/SB0/n2536 , \U1/keyexpantion/SB0/n2535 ,
         \U1/keyexpantion/SB0/n2534 , \U1/keyexpantion/SB0/n2533 ,
         \U1/keyexpantion/SB0/n2532 , \U1/keyexpantion/SB0/n2531 ,
         \U1/keyexpantion/SB0/n2530 , \U1/keyexpantion/SB0/n2529 ,
         \U1/keyexpantion/SB0/n2528 , \U1/keyexpantion/SB0/n2527 ,
         \U1/keyexpantion/SB0/n2526 , \U1/keyexpantion/SB0/n2525 ,
         \U1/keyexpantion/SB0/n2524 , \U1/keyexpantion/SB0/n2523 ,
         \U1/keyexpantion/SB0/n2522 , \U1/keyexpantion/SB0/n2521 ,
         \U1/keyexpantion/SB0/n2520 , \U1/keyexpantion/SB0/n2519 ,
         \U1/keyexpantion/SB0/n2518 , \U1/keyexpantion/SB0/n2517 ,
         \U1/keyexpantion/SB0/n2516 , \U1/keyexpantion/SB0/n2515 ,
         \U1/keyexpantion/SB0/n2514 , \U1/keyexpantion/SB0/n2513 ,
         \U1/keyexpantion/SB0/n2512 , \U1/keyexpantion/SB0/n2511 ,
         \U1/keyexpantion/SB0/n2510 , \U1/keyexpantion/SB0/n2509 ,
         \U1/keyexpantion/SB0/n2508 , \U1/keyexpantion/SB0/n2507 ,
         \U1/keyexpantion/SB0/n2506 , \U1/keyexpantion/SB0/n2505 ,
         \U1/keyexpantion/SB0/n2504 , \U1/keyexpantion/SB0/n2503 ,
         \U1/keyexpantion/SB0/n2502 , \U1/keyexpantion/SB0/n2501 ,
         \U1/keyexpantion/SB0/n2500 , \U1/keyexpantion/SB0/n2499 ,
         \U1/keyexpantion/SB0/n2498 , \U1/keyexpantion/SB0/n2497 ,
         \U1/keyexpantion/SB0/n2496 , \U1/keyexpantion/SB0/n2495 ,
         \U1/keyexpantion/SB0/n2494 , \U1/keyexpantion/SB0/n2493 ,
         \U1/keyexpantion/SB0/n2492 , \U1/keyexpantion/SB0/n2491 ,
         \U1/keyexpantion/SB0/n2490 , \U1/keyexpantion/SB0/n2489 ,
         \U1/keyexpantion/SB0/n2488 , \U1/keyexpantion/SB0/n2487 ,
         \U1/keyexpantion/SB0/n2486 , \U1/keyexpantion/SB0/n2485 ,
         \U1/keyexpantion/SB0/n2484 , \U1/keyexpantion/SB0/n2483 ,
         \U1/keyexpantion/SB0/n2482 , \U1/keyexpantion/SB0/n2481 ,
         \U1/keyexpantion/SB0/n2480 , \U1/keyexpantion/SB0/n2479 ,
         \U1/keyexpantion/SB0/n2478 , \U1/keyexpantion/SB0/n2477 ,
         \U1/keyexpantion/SB0/n2476 , \U1/keyexpantion/SB0/n2475 ,
         \U1/keyexpantion/SB0/n2474 , \U1/keyexpantion/SB0/n2473 ,
         \U1/keyexpantion/SB0/n2472 , \U1/keyexpantion/SB0/n2471 ,
         \U1/keyexpantion/SB0/n2470 , \U1/keyexpantion/SB0/n2469 ,
         \U1/keyexpantion/SB0/n2468 , \U1/keyexpantion/SB0/n2467 ,
         \U1/keyexpantion/SB0/n2466 , \U1/keyexpantion/SB0/n2465 ,
         \U1/keyexpantion/SB0/n2464 , \U1/keyexpantion/SB0/n2463 ,
         \U1/keyexpantion/SB0/n2462 , \U1/keyexpantion/SB0/n2461 ,
         \U1/keyexpantion/SB0/n2460 , \U1/keyexpantion/SB0/n2459 ,
         \U1/keyexpantion/SB0/n2458 , \U1/keyexpantion/SB0/n2457 ,
         \U1/keyexpantion/SB0/n2456 , \U1/keyexpantion/SB0/n2455 ,
         \U1/keyexpantion/SB0/n2454 , \U1/keyexpantion/SB0/n2453 ,
         \U1/keyexpantion/SB0/n2452 , \U1/keyexpantion/SB0/n2451 ,
         \U1/keyexpantion/SB0/n2450 , \U1/keyexpantion/SB0/n2449 ,
         \U1/keyexpantion/SB0/n2448 , \U1/keyexpantion/SB0/n2447 ,
         \U1/keyexpantion/SB0/n2446 , \U1/keyexpantion/SB0/n2445 ,
         \U1/keyexpantion/SB0/n2444 , \U1/keyexpantion/SB0/n2443 ,
         \U1/keyexpantion/SB0/n2442 , \U1/keyexpantion/SB0/n2441 ,
         \U1/keyexpantion/SB0/n2440 , \U1/keyexpantion/SB0/n2439 ,
         \U1/keyexpantion/SB0/n2438 , \U1/keyexpantion/SB0/n2437 ,
         \U1/keyexpantion/SB0/n2436 , \U1/keyexpantion/SB0/n2435 ,
         \U1/keyexpantion/SB0/n2434 , \U1/keyexpantion/SB0/n2433 ,
         \U1/keyexpantion/SB0/n2432 , \U1/keyexpantion/SB0/n2431 ,
         \U1/keyexpantion/SB0/n2430 , \U1/keyexpantion/SB0/n2429 ,
         \U1/keyexpantion/SB0/n2428 , \U1/keyexpantion/SB0/n2427 ,
         \U1/keyexpantion/SB0/n2426 , \U1/keyexpantion/SB0/n2425 ,
         \U1/keyexpantion/SB0/n2424 , \U1/keyexpantion/SB0/n2423 ,
         \U1/keyexpantion/SB0/n2422 , \U1/keyexpantion/SB0/n2421 ,
         \U1/keyexpantion/SB0/n2420 , \U1/keyexpantion/SB0/n2419 ,
         \U1/keyexpantion/SB0/n2418 , \U1/keyexpantion/SB0/n2417 ,
         \U1/keyexpantion/SB0/n2416 , \U1/keyexpantion/SB0/n2415 ,
         \U1/keyexpantion/SB0/n2414 , \U1/keyexpantion/SB0/n2413 ,
         \U1/keyexpantion/SB0/n2412 , \U1/keyexpantion/SB0/n2411 ,
         \U1/keyexpantion/SB0/n2410 , \U1/keyexpantion/SB0/n2409 ,
         \U1/keyexpantion/SB0/n2408 , \U1/keyexpantion/SB0/n2407 ,
         \U1/keyexpantion/SB0/n2406 , \U1/keyexpantion/SB0/n2405 ,
         \U1/keyexpantion/SB0/n2404 , \U1/keyexpantion/SB0/n2403 ,
         \U1/keyexpantion/SB0/n2402 , \U1/keyexpantion/SB0/n2401 ,
         \U1/keyexpantion/SB0/n2400 , \U1/keyexpantion/SB0/n2399 ,
         \U1/keyexpantion/SB0/n2398 , \U1/keyexpantion/SB0/n2397 ,
         \U1/keyexpantion/SB0/n2396 , \U1/keyexpantion/SB0/n2395 ,
         \U1/keyexpantion/SB0/n2394 , \U1/keyexpantion/SB0/n2393 ,
         \U1/keyexpantion/SB0/n2392 , \U1/keyexpantion/SB0/n2391 ,
         \U1/keyexpantion/SB0/n2390 , \U1/keyexpantion/SB0/n2389 ,
         \U1/keyexpantion/SB0/n2388 , \U1/keyexpantion/SB0/n2387 ,
         \U1/keyexpantion/SB0/n2386 , \U1/keyexpantion/SB0/n2385 ,
         \U1/keyexpantion/SB0/n2384 , \U1/keyexpantion/SB0/n2383 ,
         \U1/keyexpantion/SB0/n2382 , \U1/keyexpantion/SB0/n2381 ,
         \U1/keyexpantion/SB0/n2380 , \U1/keyexpantion/SB0/n2379 ,
         \U1/keyexpantion/SB0/n2378 , \U1/keyexpantion/SB0/n2377 ,
         \U1/keyexpantion/SB0/n2376 , \U1/keyexpantion/SB0/n2375 ,
         \U1/keyexpantion/SB0/n2374 , \U1/keyexpantion/SB0/n2373 ,
         \U1/keyexpantion/SB0/n2372 , \U1/keyexpantion/SB0/n2371 ,
         \U1/keyexpantion/SB0/n2370 , \U1/keyexpantion/SB0/n2369 ,
         \U1/keyexpantion/SB0/n2368 , \U1/keyexpantion/SB0/n2367 ,
         \U1/keyexpantion/SB0/n2366 , \U1/keyexpantion/SB0/n2365 ,
         \U1/keyexpantion/SB0/n2364 , \U1/keyexpantion/SB0/n2363 ,
         \U1/keyexpantion/SB0/n2362 , \U1/keyexpantion/SB0/n2361 ,
         \U1/keyexpantion/SB0/n2360 , \U1/keyexpantion/SB0/n2359 ,
         \U1/keyexpantion/SB0/n2358 , \U1/keyexpantion/SB0/n2357 ,
         \U1/keyexpantion/SB0/n2356 , \U1/keyexpantion/SB0/n2355 ,
         \U1/keyexpantion/SB0/n2354 , \U1/keyexpantion/SB0/n2353 ,
         \U1/keyexpantion/SB0/n2352 , \U1/keyexpantion/SB0/n2351 ,
         \U1/keyexpantion/SB0/n2350 , \U1/keyexpantion/SB0/n2349 ,
         \U1/keyexpantion/SB0/n2348 , \U1/keyexpantion/SB0/n2347 ,
         \U1/keyexpantion/SB0/n2346 , \U1/keyexpantion/SB0/n2345 ,
         \U1/keyexpantion/SB0/n2344 , \U1/keyexpantion/SB0/n2343 ,
         \U1/keyexpantion/SB0/n2342 , \U1/keyexpantion/SB0/n2341 ,
         \U1/keyexpantion/SB0/n2340 , \U1/keyexpantion/SB0/n2339 ,
         \U1/keyexpantion/SB0/n2338 , \U1/keyexpantion/SB0/n2337 ,
         \U1/keyexpantion/SB0/n2336 , \U1/keyexpantion/SB0/n2335 ,
         \U1/keyexpantion/SB0/n2334 , \U1/keyexpantion/SB0/n2333 ,
         \U1/keyexpantion/SB0/n2332 , \U1/keyexpantion/SB0/n2331 ,
         \U1/keyexpantion/SB0/n2330 , \U1/keyexpantion/SB0/n2329 ,
         \U1/keyexpantion/SB0/n2328 , \U1/keyexpantion/SB0/n2327 ,
         \U1/keyexpantion/SB0/n2326 , \U1/keyexpantion/SB0/n2325 ,
         \U1/keyexpantion/SB0/n2324 , \U1/keyexpantion/SB0/n2323 ,
         \U1/keyexpantion/SB0/n2322 , \U1/keyexpantion/SB0/n2321 ,
         \U1/keyexpantion/SB0/n2320 , \U1/keyexpantion/SB0/n2319 ,
         \U1/keyexpantion/SB0/n2318 , \U1/keyexpantion/SB0/n2317 ,
         \U1/keyexpantion/SB0/n2316 , \U1/keyexpantion/SB0/n2315 ,
         \U1/keyexpantion/SB0/n2314 , \U1/keyexpantion/SB0/n2313 ,
         \U1/keyexpantion/SB0/n2312 , \U1/keyexpantion/SB0/n2311 ,
         \U1/keyexpantion/SB0/n2310 , \U1/keyexpantion/SB0/n2309 ,
         \U1/keyexpantion/SB0/n2308 , \U1/keyexpantion/SB0/n2307 ,
         \U1/keyexpantion/SB0/n2306 , \U1/keyexpantion/SB0/n2305 ,
         \U1/keyexpantion/SB0/n2304 , \U1/keyexpantion/SB0/n2303 ,
         \U1/keyexpantion/SB0/n2302 , \U1/keyexpantion/SB0/n2301 ,
         \U1/keyexpantion/SB0/n2300 , \U1/keyexpantion/SB0/n2299 ,
         \U1/keyexpantion/SB0/n2298 , \U1/keyexpantion/SB0/n2297 ,
         \U1/keyexpantion/SB0/n2296 , \U1/keyexpantion/SB0/n2295 ,
         \U1/keyexpantion/SB0/n2294 , \U1/keyexpantion/SB0/n2293 ,
         \U1/keyexpantion/SB0/n2292 , \U1/keyexpantion/SB0/n2291 ,
         \U1/keyexpantion/SB0/n2290 , \U1/keyexpantion/SB0/n2289 ,
         \U1/keyexpantion/SB0/n2288 , \U1/keyexpantion/SB0/n2287 ,
         \U1/keyexpantion/SB0/n2286 , \U1/keyexpantion/SB0/n2285 ,
         \U1/keyexpantion/SB0/n2284 , \U1/keyexpantion/SB0/n2283 ,
         \U1/keyexpantion/SB0/n2282 , \U1/keyexpantion/SB0/n2281 ,
         \U1/keyexpantion/SB0/n2280 , \U1/keyexpantion/SB0/n2279 ,
         \U1/keyexpantion/SB0/n2278 , \U1/keyexpantion/SB0/n2277 ,
         \U1/keyexpantion/SB0/n2276 , \U1/keyexpantion/SB0/n2275 ,
         \U1/keyexpantion/SB0/n2274 , \U1/keyexpantion/SB0/n2273 ,
         \U1/keyexpantion/SB0/n2272 , \U1/keyexpantion/SB0/n2271 ,
         \U1/keyexpantion/SB0/n2270 , \U1/keyexpantion/SB0/n2269 ,
         \U1/keyexpantion/SB0/n2268 , \U1/keyexpantion/SB0/n2267 ,
         \U1/keyexpantion/SB0/n2266 , \U1/keyexpantion/SB0/n2265 ,
         \U1/keyexpantion/SB0/n2264 , \U1/keyexpantion/SB0/n2263 ,
         \U1/keyexpantion/SB0/n2262 , \U1/keyexpantion/SB0/n2261 ,
         \U1/keyexpantion/SB0/n2260 , \U1/keyexpantion/SB0/n2259 ,
         \U1/keyexpantion/SB0/n2258 , \U1/keyexpantion/SB0/n2257 ,
         \U1/keyexpantion/SB0/n2256 , \U1/keyexpantion/SB0/n2255 ,
         \U1/keyexpantion/SB0/n2254 , \U1/keyexpantion/SB0/n2253 ,
         \U1/keyexpantion/SB0/n2252 , \U1/keyexpantion/SB0/n2251 ,
         \U1/keyexpantion/SB0/n2250 , \U1/keyexpantion/SB0/n2249 ,
         \U1/keyexpantion/SB0/n2248 , \U1/keyexpantion/SB0/n2247 ,
         \U1/keyexpantion/SB0/n2246 , \U1/keyexpantion/SB0/n2245 ,
         \U1/keyexpantion/SB0/n2244 , \U1/keyexpantion/SB0/n2243 ,
         \U1/keyexpantion/SB0/n2242 , \U1/keyexpantion/SB0/n2241 ,
         \U1/keyexpantion/SB0/n2240 , \U1/keyexpantion/SB0/n2239 ,
         \U1/keyexpantion/SB0/n2238 , \U1/keyexpantion/SB0/n2237 ,
         \U1/keyexpantion/SB0/n2236 , \U1/keyexpantion/SB0/n2235 ,
         \U1/keyexpantion/SB0/n2234 , \U1/keyexpantion/SB0/n2233 ,
         \U1/keyexpantion/SB0/n2232 , \U1/keyexpantion/SB0/n2231 ,
         \U1/keyexpantion/SB0/n2230 , \U1/keyexpantion/SB0/n2229 ,
         \U1/keyexpantion/SB0/n2228 , \U1/keyexpantion/SB0/n2227 ,
         \U1/keyexpantion/SB0/n2226 , \U1/keyexpantion/SB0/n2225 ,
         \U1/keyexpantion/SB0/n2224 , \U1/keyexpantion/SB0/n2223 ,
         \U1/keyexpantion/SB0/n2222 , \U1/keyexpantion/SB0/n2221 ,
         \U1/keyexpantion/SB0/n2220 , \U1/keyexpantion/SB0/n2219 ,
         \U1/keyexpantion/SB0/n2218 , \U1/keyexpantion/SB0/n2217 ,
         \U1/keyexpantion/SB0/n2216 , \U1/keyexpantion/SB0/n2215 ,
         \U1/keyexpantion/SB0/n2214 , \U1/keyexpantion/SB0/n2213 ,
         \U1/keyexpantion/SB0/n2212 , \U1/keyexpantion/SB0/n2211 ,
         \U1/keyexpantion/SB0/n2210 , \U1/keyexpantion/SB0/n2209 ,
         \U1/keyexpantion/SB0/n2208 , \U1/keyexpantion/SB0/n2207 ,
         \U1/keyexpantion/SB0/n2206 , \U1/keyexpantion/SB0/n2205 ,
         \U1/keyexpantion/SB0/n2204 , \U1/keyexpantion/SB0/n2203 ,
         \U1/keyexpantion/SB0/n2202 , \U1/keyexpantion/SB0/n2201 ,
         \U1/keyexpantion/SB0/n2200 , \U1/keyexpantion/SB0/n2199 ,
         \U1/keyexpantion/SB0/n2198 , \U1/keyexpantion/SB0/n2197 ,
         \U1/keyexpantion/SB0/n2196 , \U1/keyexpantion/SB0/n2195 ,
         \U1/keyexpantion/SB0/n2194 , \U1/keyexpantion/SB0/n2193 ,
         \U1/keyexpantion/SB0/n2192 , \U1/keyexpantion/SB0/n2191 ,
         \U1/keyexpantion/SB0/n2190 , \U1/keyexpantion/SB0/n2189 ,
         \U1/keyexpantion/SB0/n2188 , \U1/keyexpantion/SB0/n2187 ,
         \U1/keyexpantion/SB0/n2186 , \U1/keyexpantion/SB0/n2185 ,
         \U1/keyexpantion/SB0/n2184 , \U1/keyexpantion/SB0/n2183 ,
         \U1/keyexpantion/SB0/n2182 , \U1/keyexpantion/SB0/n2181 ,
         \U1/keyexpantion/SB0/n2180 , \U1/keyexpantion/SB0/n2179 ,
         \U1/keyexpantion/SB0/n2178 , \U1/keyexpantion/SB0/n2177 ,
         \U1/keyexpantion/SB0/n2176 , \U1/keyexpantion/SB0/n2175 ,
         \U1/keyexpantion/SB0/n2174 , \U1/keyexpantion/SB0/n2173 ,
         \U1/keyexpantion/SB0/n2172 , \U1/keyexpantion/SB0/n2171 ,
         \U1/keyexpantion/SB0/n2170 , \U1/keyexpantion/SB0/n2169 ,
         \U1/keyexpantion/SB0/n2168 , \U1/keyexpantion/SB0/n2167 ,
         \U1/keyexpantion/SB0/n2166 , \U1/keyexpantion/SB0/n2165 ,
         \U1/keyexpantion/SB0/n2164 , \U1/keyexpantion/SB0/n2163 ,
         \U1/keyexpantion/SB0/n2162 , \U1/keyexpantion/SB0/n2161 ,
         \U1/keyexpantion/SB0/n2160 , \U1/keyexpantion/SB0/n2159 ,
         \U1/keyexpantion/SB0/n2158 , \U1/keyexpantion/SB0/n2157 ,
         \U1/keyexpantion/SB0/n2156 , \U1/keyexpantion/SB0/n2155 ,
         \U1/keyexpantion/SB0/n2154 , \U1/keyexpantion/SB0/n2153 ,
         \U1/keyexpantion/SB0/n2152 , \U1/keyexpantion/SB0/n2151 ,
         \U1/keyexpantion/SB0/n2150 , \U1/keyexpantion/SB0/n2149 ,
         \U1/keyexpantion/SB0/n2148 , \U1/keyexpantion/SB0/n2147 ,
         \U1/keyexpantion/SB0/n2146 , \U1/keyexpantion/SB0/n2145 ,
         \U1/keyexpantion/SB0/n2144 , \U1/keyexpantion/SB0/n2143 ,
         \U1/keyexpantion/SB0/n2142 , \U1/keyexpantion/SB0/n2141 ,
         \U1/keyexpantion/SB0/n2140 , \U1/keyexpantion/SB0/n2139 ,
         \U1/keyexpantion/SB0/n2138 , \U1/keyexpantion/SB0/n2137 ,
         \U1/keyexpantion/SB0/n2136 , \U1/keyexpantion/SB0/n2135 ,
         \U1/keyexpantion/SB0/n2134 , \U1/keyexpantion/SB0/n2133 ,
         \U1/keyexpantion/SB0/n2132 , \U1/keyexpantion/SB0/n2131 ,
         \U1/keyexpantion/SB0/n2130 , \U1/keyexpantion/SB0/n2129 ,
         \U1/keyexpantion/SB0/n2128 , \U1/keyexpantion/SB0/n2127 ,
         \U1/keyexpantion/SB0/n2126 , \U1/keyexpantion/SB0/n2125 ,
         \U1/keyexpantion/SB0/n2124 , \U1/keyexpantion/SB0/n2123 ,
         \U1/keyexpantion/SB0/n2122 , \U1/keyexpantion/SB0/n2121 ,
         \U1/keyexpantion/SB0/n2120 , \U1/keyexpantion/SB0/n2119 ,
         \U1/keyexpantion/SB0/n2118 , \U1/keyexpantion/SB0/n2117 ,
         \U1/keyexpantion/SB0/n2116 , \U1/keyexpantion/SB0/n2115 ,
         \U1/keyexpantion/SB0/n2114 , \U1/keyexpantion/SB0/n2113 ,
         \U1/keyexpantion/SB0/n2112 , \U1/keyexpantion/SB0/n2111 ,
         \U1/keyexpantion/SB0/n2110 , \U1/keyexpantion/SB0/n2109 ,
         \U1/keyexpantion/SB0/n2108 , \U1/keyexpantion/SB0/n2107 ,
         \U1/keyexpantion/SB0/n2106 , \U1/keyexpantion/SB0/n2105 ,
         \U1/keyexpantion/SB0/n2104 , \U1/keyexpantion/SB0/n2103 ,
         \U1/keyexpantion/SB0/n2102 , \U1/keyexpantion/SB0/n2101 ,
         \U1/keyexpantion/SB0/n2100 , \U1/keyexpantion/SB0/n2099 ,
         \U1/keyexpantion/SB0/n2098 , \U1/keyexpantion/SB0/n2097 ,
         \U1/keyexpantion/SB0/n2096 , \U1/keyexpantion/SB0/n2095 ,
         \U1/keyexpantion/SB0/n2094 , \U1/keyexpantion/SB0/n2093 ,
         \U1/keyexpantion/SB0/n2092 , \U1/keyexpantion/SB0/n2091 ,
         \U1/keyexpantion/SB0/n2090 , \U1/keyexpantion/SB0/n2089 ,
         \U1/keyexpantion/SB0/n2088 , \U1/keyexpantion/SB0/n2087 ,
         \U1/keyexpantion/SB0/n2086 , \U1/keyexpantion/SB0/n2085 ,
         \U1/keyexpantion/SB0/n2084 , \U1/keyexpantion/SB0/n2083 ,
         \U1/keyexpantion/SB0/n2082 , \U1/keyexpantion/SB0/n2081 ,
         \U1/keyexpantion/SB0/n2080 , \U1/keyexpantion/SB0/n2079 ,
         \U1/keyexpantion/SB0/n2078 , \U1/keyexpantion/SB0/n2077 ,
         \U1/keyexpantion/SB0/n2076 , \U1/keyexpantion/SB0/n2075 ,
         \U1/keyexpantion/SB0/n2074 , \U1/keyexpantion/SB0/n2073 ,
         \U1/keyexpantion/SB0/n2072 , \U1/keyexpantion/SB0/n2071 ,
         \U1/keyexpantion/SB0/n2070 , \U1/keyexpantion/SB0/n2069 ,
         \U1/keyexpantion/SB0/n2068 , \U1/keyexpantion/SB0/n2067 ,
         \U1/keyexpantion/SB0/n2066 , \U1/keyexpantion/SB0/n2065 ,
         \U1/keyexpantion/SB0/n2064 , \U1/keyexpantion/SB0/n2063 ,
         \U1/keyexpantion/SB0/n2062 , \U1/keyexpantion/SB0/n2061 ,
         \U1/keyexpantion/SB0/n2060 , \U1/keyexpantion/SB0/n2059 ,
         \U1/keyexpantion/SB0/n2058 , \U1/keyexpantion/SB0/n2057 ,
         \U1/keyexpantion/SB0/n2056 , \U1/keyexpantion/SB0/n2055 ,
         \U1/keyexpantion/SB0/n2054 , \U1/keyexpantion/SB0/n2053 ,
         \U1/keyexpantion/SB0/n2052 , \U1/keyexpantion/SB0/n2051 ,
         \U1/keyexpantion/SB0/n2050 , \U1/keyexpantion/SB0/n2049 ,
         \U1/keyexpantion/SB0/n2048 , \U1/keyexpantion/SB0/n2047 ,
         \U1/keyexpantion/SB0/n2046 , \U1/keyexpantion/SB0/n2045 ,
         \U1/keyexpantion/SB0/n2044 , \U1/keyexpantion/SB0/n2043 ,
         \U1/keyexpantion/SB0/n2042 , \U1/keyexpantion/SB0/n2041 ,
         \U1/keyexpantion/SB0/n2040 , \U1/keyexpantion/SB0/n2039 ,
         \U1/keyexpantion/SB0/n2038 , \U1/keyexpantion/SB0/n2037 ,
         \U1/keyexpantion/SB0/n2036 , \U1/keyexpantion/SB0/n2035 ,
         \U1/keyexpantion/SB0/n2034 , \U1/keyexpantion/SB0/n2033 ,
         \U1/keyexpantion/SB0/n2032 , \U1/keyexpantion/SB0/n2031 ,
         \U1/keyexpantion/SB0/n2030 , \U1/keyexpantion/SB0/n2029 ,
         \U1/keyexpantion/SB0/n2028 , \U1/keyexpantion/SB0/n2027 ,
         \U1/keyexpantion/SB0/n2026 , \U1/keyexpantion/SB0/n2025 ,
         \U1/keyexpantion/SB0/n2024 , \U1/keyexpantion/SB0/n2023 ,
         \U1/keyexpantion/SB0/n2022 , \U1/keyexpantion/SB0/n2021 ,
         \U1/keyexpantion/SB0/n2020 , \U1/keyexpantion/SB0/n2019 ,
         \U1/keyexpantion/SB0/n2018 , \U1/keyexpantion/SB0/n2017 ,
         \U1/keyexpantion/SB0/n2016 , \U1/keyexpantion/SB0/n2015 ,
         \U1/keyexpantion/SB0/n2014 , \U1/keyexpantion/SB0/n2013 ,
         \U1/keyexpantion/SB0/n2012 , \U1/keyexpantion/SB0/n2011 ,
         \U1/keyexpantion/SB0/n2010 , \U1/keyexpantion/SB0/n2009 ,
         \U1/keyexpantion/SB0/n2008 , \U1/keyexpantion/SB0/n2007 ,
         \U1/keyexpantion/SB0/n2006 , \U1/keyexpantion/SB0/n2005 ,
         \U1/keyexpantion/SB0/n2004 , \U1/keyexpantion/SB0/n2003 ,
         \U1/keyexpantion/SB0/n2002 , \U1/keyexpantion/SB0/n2001 ,
         \U1/keyexpantion/SB0/n2000 , \U1/keyexpantion/SB0/n1999 ,
         \U1/keyexpantion/SB0/n1998 , \U1/keyexpantion/SB0/n1997 ,
         \U1/keyexpantion/SB0/n1996 , \U1/keyexpantion/SB0/n1995 ,
         \U1/keyexpantion/SB0/n1994 , \U1/keyexpantion/SB0/n1993 ,
         \U1/keyexpantion/SB0/n1992 , \U1/keyexpantion/SB0/n1991 ,
         \U1/keyexpantion/SB0/n1990 , \U1/keyexpantion/SB0/n1989 ,
         \U1/keyexpantion/SB0/n1988 , \U1/keyexpantion/SB0/n1987 ,
         \U1/keyexpantion/SB0/n1986 , \U1/keyexpantion/SB0/n1985 ,
         \U1/keyexpantion/SB0/n1984 , \U1/keyexpantion/SB0/n1983 ,
         \U1/keyexpantion/SB0/n1982 , \U1/keyexpantion/SB0/n1981 ,
         \U1/keyexpantion/SB0/n1980 , \U1/keyexpantion/SB0/n1979 ,
         \U1/keyexpantion/SB0/n1978 , \U1/keyexpantion/SB0/n1977 ,
         \U1/keyexpantion/SB0/n1976 , \U1/keyexpantion/SB0/n1975 ,
         \U1/keyexpantion/SB0/n1974 , \U1/keyexpantion/SB0/n1973 ,
         \U1/keyexpantion/SB0/n1972 , \U1/keyexpantion/SB0/n1971 ,
         \U1/keyexpantion/SB0/n1970 , \U1/keyexpantion/SB0/n1969 ,
         \U1/keyexpantion/SB0/n1968 , \U1/keyexpantion/SB0/n1967 ,
         \U1/keyexpantion/SB0/n1966 , \U1/keyexpantion/SB0/n1965 ,
         \U1/keyexpantion/SB0/n1964 , \U1/keyexpantion/SB0/n1963 ,
         \U1/keyexpantion/SB0/n1962 , \U1/keyexpantion/SB0/n1961 ,
         \U1/keyexpantion/SB0/n1960 , \U1/keyexpantion/SB0/n1959 ,
         \U1/keyexpantion/SB0/n1958 , \U1/keyexpantion/SB0/n1957 ,
         \U1/keyexpantion/SB0/n1956 , \U1/keyexpantion/SB0/n1955 ,
         \U1/keyexpantion/SB0/n1954 , \U1/keyexpantion/SB0/n1953 ,
         \U1/keyexpantion/SB0/n1952 , \U1/keyexpantion/SB0/n1951 ,
         \U1/keyexpantion/SB0/n1950 , \U1/keyexpantion/SB0/n1949 ,
         \U1/keyexpantion/SB0/n1948 , \U1/keyexpantion/SB0/n1947 ,
         \U1/keyexpantion/SB0/n1946 , \U1/keyexpantion/SB0/n1945 ,
         \U1/keyexpantion/SB0/n1944 , \U1/keyexpantion/SB0/n1943 ,
         \U1/keyexpantion/SB0/n1942 , \U1/keyexpantion/SB0/n1941 ,
         \U1/keyexpantion/SB0/n1940 , \U1/keyexpantion/SB0/n1939 ,
         \U1/keyexpantion/SB0/n1938 , \U1/keyexpantion/SB0/n1937 ,
         \U1/keyexpantion/SB0/n1936 , \U1/keyexpantion/SB0/n1935 ,
         \U1/keyexpantion/SB0/n1934 , \U1/keyexpantion/SB0/n1933 ,
         \U1/keyexpantion/SB0/n1932 , \U1/keyexpantion/SB0/n1931 ,
         \U1/keyexpantion/SB0/n1930 , \U1/keyexpantion/SB0/n1929 ,
         \U1/keyexpantion/SB0/n1928 , \U1/keyexpantion/SB0/n1927 ,
         \U1/keyexpantion/SB0/n1926 , \U1/keyexpantion/SB0/n1925 ,
         \U1/keyexpantion/SB0/n1924 , \U1/keyexpantion/SB0/n1923 ,
         \U1/keyexpantion/SB0/n1922 , \U1/keyexpantion/SB0/n1921 ,
         \U1/keyexpantion/SB0/n1920 , \U1/keyexpantion/SB0/n1919 ,
         \U1/keyexpantion/SB0/n1918 , \U1/keyexpantion/SB0/n1917 ,
         \U1/keyexpantion/SB0/n1916 , \U1/keyexpantion/SB0/n1915 ,
         \U1/keyexpantion/SB0/n1914 , \U1/keyexpantion/SB0/n1913 ,
         \U1/keyexpantion/SB0/n1912 , \U1/keyexpantion/SB0/n1911 ,
         \U1/keyexpantion/SB0/n1910 , \U1/keyexpantion/SB0/n1909 ,
         \U1/keyexpantion/SB0/n1908 , \U1/keyexpantion/SB0/n1907 ,
         \U1/keyexpantion/SB0/n1906 , \U1/keyexpantion/SB0/n1905 ,
         \U1/keyexpantion/SB0/n1904 , \U1/keyexpantion/SB0/n1903 ,
         \U1/keyexpantion/SB0/n1902 , \U1/keyexpantion/SB0/n1901 ,
         \U1/keyexpantion/SB0/n1900 , \U1/keyexpantion/SB0/n1899 ,
         \U1/keyexpantion/SB0/n1898 , \U1/keyexpantion/SB0/n1897 ,
         \U1/keyexpantion/SB0/n1896 , \U1/keyexpantion/SB0/n1895 ,
         \U1/keyexpantion/SB0/n1894 , \U1/keyexpantion/SB0/n1893 ,
         \U1/keyexpantion/SB0/n1892 , \U1/keyexpantion/SB0/n1891 ,
         \U1/keyexpantion/SB0/n1890 , \U1/keyexpantion/SB0/n1889 ,
         \U1/keyexpantion/SB0/n1888 , \U1/keyexpantion/SB0/n1887 ,
         \U1/keyexpantion/SB0/n1886 , \U1/keyexpantion/SB0/n1885 ,
         \U1/keyexpantion/SB0/n1884 , \U1/keyexpantion/SB0/n1883 ,
         \U1/keyexpantion/SB0/n1882 , \U1/keyexpantion/SB0/n1881 ,
         \U1/keyexpantion/SB0/n1880 , \U1/keyexpantion/SB0/n1879 ,
         \U1/keyexpantion/SB0/n1878 , \U1/keyexpantion/SB0/n1877 ,
         \U1/keyexpantion/SB0/n1876 , \U1/keyexpantion/SB0/n1875 ,
         \U1/keyexpantion/SB0/n1874 , \U1/keyexpantion/SB0/n1873 ,
         \U1/keyexpantion/SB0/n1872 , \U1/keyexpantion/SB0/n1871 ,
         \U1/keyexpantion/SB0/n1870 , \U1/keyexpantion/SB0/n1869 ,
         \U1/keyexpantion/SB0/n1868 , \U1/keyexpantion/SB0/n1867 ,
         \U1/keyexpantion/SB0/n1866 , \U1/keyexpantion/SB0/n1865 ,
         \U1/keyexpantion/SB0/n1864 , \U1/keyexpantion/SB0/n1863 ,
         \U1/keyexpantion/SB0/n1862 , \U1/keyexpantion/SB0/n1861 ,
         \U1/keyexpantion/SB0/n1860 , \U1/keyexpantion/SB0/n1859 ,
         \U1/keyexpantion/SB0/n1858 , \U1/keyexpantion/SB0/n1857 ,
         \U1/keyexpantion/SB0/n1856 , \U1/keyexpantion/SB0/n1855 ,
         \U1/keyexpantion/SB0/n1854 , \U1/keyexpantion/SB0/n1853 ,
         \U1/keyexpantion/SB0/n1852 , \U1/keyexpantion/SB0/n1851 ,
         \U1/keyexpantion/SB0/n1850 , \U1/keyexpantion/SB0/n1849 ,
         \U1/keyexpantion/SB0/n1848 , \U1/keyexpantion/SB0/n1847 ,
         \U1/keyexpantion/SB0/n1846 , \U1/keyexpantion/SB0/n1845 ,
         \U1/keyexpantion/SB0/n1844 , \U1/keyexpantion/SB0/n1843 ,
         \U1/keyexpantion/SB0/n1842 , \U1/keyexpantion/SB0/n1841 ,
         \U1/keyexpantion/SB0/n1840 , \U1/keyexpantion/SB0/n1839 ,
         \U1/keyexpantion/SB0/n1838 , \U1/keyexpantion/SB0/n1837 ,
         \U1/keyexpantion/SB0/n1836 , \U1/keyexpantion/SB0/n1835 ,
         \U1/keyexpantion/SB0/n1834 , \U1/keyexpantion/SB0/n1833 ,
         \U1/keyexpantion/SB0/n1832 , \U1/keyexpantion/SB0/n1831 ,
         \U1/keyexpantion/SB0/n1830 , \U1/keyexpantion/SB0/n1829 ,
         \U1/keyexpantion/SB0/n1828 , \U1/keyexpantion/SB0/n1827 ,
         \U1/keyexpantion/SB0/n1826 , \U1/keyexpantion/SB0/n1825 ,
         \U1/keyexpantion/SB0/n1824 , \U1/keyexpantion/SB0/n1823 ,
         \U1/keyexpantion/SB0/n1822 , \U1/keyexpantion/SB0/n1821 ,
         \U1/keyexpantion/SB0/n1820 , \U1/keyexpantion/SB0/n1819 ,
         \U1/keyexpantion/SB0/n1818 , \U1/keyexpantion/SB0/n1817 ,
         \U1/keyexpantion/SB0/n1816 , \U1/keyexpantion/SB0/n1815 ,
         \U1/keyexpantion/SB0/n1814 , \U1/keyexpantion/SB0/n1813 ,
         \U1/keyexpantion/SB0/n1812 , \U1/keyexpantion/SB0/n1811 ,
         \U1/keyexpantion/SB0/n1810 , \U1/keyexpantion/SB0/n1809 ,
         \U1/keyexpantion/SB0/n1808 , \U1/keyexpantion/SB0/n1807 ,
         \U1/keyexpantion/SB0/n1806 , \U1/keyexpantion/SB0/n1805 ,
         \U1/keyexpantion/SB0/n1804 , \U1/keyexpantion/SB0/n1803 ,
         \U1/keyexpantion/SB0/n1802 , \U1/keyexpantion/SB0/n1801 ,
         \U1/keyexpantion/SB0/n1800 , \U1/keyexpantion/SB0/n1799 ,
         \U1/keyexpantion/SB0/n1798 , \U1/keyexpantion/SB0/n1797 ,
         \U1/keyexpantion/SB0/n1796 , \U1/keyexpantion/SB0/n1795 ,
         \U1/keyexpantion/SB0/n1794 , \U1/keyexpantion/SB0/n1793 ,
         \U1/keyexpantion/SB0/n1792 , \U1/keyexpantion/SB0/n1791 ,
         \U1/keyexpantion/SB0/n1790 , \U1/keyexpantion/SB0/n1789 ,
         \U1/keyexpantion/SB0/n1788 , \U1/keyexpantion/SB0/n1787 ,
         \U1/keyexpantion/SB0/n1786 , \U1/keyexpantion/SB0/n1785 ,
         \U1/keyexpantion/SB0/n1784 , \U1/keyexpantion/SB0/n1783 ,
         \U1/keyexpantion/SB0/n1782 , \U1/keyexpantion/SB0/n1781 ,
         \U1/keyexpantion/SB0/n1780 , \U1/keyexpantion/SB0/n1779 ,
         \U1/keyexpantion/SB0/n1778 , \U1/keyexpantion/SB0/n1777 ,
         \U1/keyexpantion/SB0/n1776 , \U1/keyexpantion/SB0/n1775 ,
         \U1/keyexpantion/SB0/n1774 , \U1/keyexpantion/SB0/n1773 ,
         \U1/keyexpantion/SB0/n1772 , \U1/keyexpantion/SB0/n1771 ,
         \U1/keyexpantion/SB0/n1770 , \U1/keyexpantion/SB0/n1769 ,
         \U1/keyexpantion/SB0/n1768 , \U1/keyexpantion/SB0/n1767 ,
         \U1/keyexpantion/SB0/n1766 , \U1/keyexpantion/SB0/n1765 ,
         \U1/keyexpantion/SB0/n1764 , \U1/keyexpantion/SB0/n1763 ,
         \U1/keyexpantion/SB0/n1762 , \U1/keyexpantion/SB0/n1761 ,
         \U1/keyexpantion/SB0/n1760 , \U1/keyexpantion/SB0/n1759 ,
         \U1/keyexpantion/SB0/n1758 , \U1/keyexpantion/SB0/n1757 ,
         \U1/keyexpantion/SB0/n1756 , \U1/keyexpantion/SB0/n1755 ,
         \U1/keyexpantion/SB0/n1754 , \U1/keyexpantion/SB0/n1753 ,
         \U1/keyexpantion/SB0/n1752 , \U1/keyexpantion/SB0/n1751 ,
         \U1/keyexpantion/SB0/n1750 , \U1/keyexpantion/SB0/n1749 ,
         \U1/keyexpantion/SB0/n1748 , \U1/keyexpantion/SB0/n1747 ,
         \U1/keyexpantion/SB0/n1746 , \U1/keyexpantion/SB0/n1745 ,
         \U1/keyexpantion/SB0/n1744 , \U1/keyexpantion/SB0/n1743 ,
         \U1/keyexpantion/SB0/n1742 , \U1/keyexpantion/SB0/n1741 ,
         \U1/keyexpantion/SB0/n1740 , \U1/keyexpantion/SB0/n1739 ,
         \U1/keyexpantion/SB0/n1738 , \U1/keyexpantion/SB0/n1737 ,
         \U1/keyexpantion/SB0/n1736 , \U1/keyexpantion/SB0/n1735 ,
         \U1/keyexpantion/SB0/n1734 , \U1/keyexpantion/SB0/n1733 ,
         \U1/keyexpantion/SB0/n1732 , \U1/keyexpantion/SB0/n1731 ,
         \U1/keyexpantion/SB0/n1730 , \U1/keyexpantion/SB0/n1729 ,
         \U1/keyexpantion/SB0/n1728 , \U1/keyexpantion/SB0/n1727 ,
         \U1/keyexpantion/SB0/n1726 , \U1/keyexpantion/SB0/n1725 ,
         \U1/keyexpantion/SB0/n1724 , \U1/keyexpantion/SB0/n1723 ,
         \U1/keyexpantion/SB0/n1722 , \U1/keyexpantion/SB0/n1721 ,
         \U1/keyexpantion/SB0/n1720 , \U1/keyexpantion/SB0/n1719 ,
         \U1/keyexpantion/SB0/n1718 , \U1/keyexpantion/SB0/n1717 ,
         \U1/keyexpantion/SB0/n1716 , \U1/keyexpantion/SB0/n1715 ,
         \U1/keyexpantion/SB0/n1714 , \U1/keyexpantion/SB0/n1713 ,
         \U1/keyexpantion/SB0/n1712 , \U1/keyexpantion/SB0/n1711 ,
         \U1/keyexpantion/SB0/n1710 , \U1/keyexpantion/SB0/n1709 ,
         \U1/keyexpantion/SB0/n1708 , \U1/keyexpantion/SB0/n1707 ,
         \U1/keyexpantion/SB0/n1706 , \U1/keyexpantion/SB0/n1705 ,
         \U1/keyexpantion/SB0/n1704 , \U1/keyexpantion/SB0/n1703 ,
         \U1/keyexpantion/SB0/n1702 , \U1/keyexpantion/SB0/n1701 ,
         \U1/keyexpantion/SB0/n1700 , \U1/keyexpantion/SB0/n1699 ,
         \U1/keyexpantion/SB0/n1698 , \U1/keyexpantion/SB0/n1697 ,
         \U1/keyexpantion/SB0/n1696 , \U1/keyexpantion/SB0/n1695 ,
         \U1/keyexpantion/SB0/n1694 , \U1/keyexpantion/SB0/n1693 ,
         \U1/keyexpantion/SB0/n1692 , \U1/keyexpantion/SB0/n1691 ,
         \U1/keyexpantion/SB0/n1690 , \U1/keyexpantion/SB0/n1689 ,
         \U1/keyexpantion/SB0/n1688 , \U1/keyexpantion/SB0/n1687 ,
         \U1/keyexpantion/SB0/n1686 , \U1/keyexpantion/SB0/n1685 ,
         \U1/keyexpantion/SB0/n1203 , \U1/keyexpantion/SB0/n1158 ,
         \U1/keyexpantion/SB0/n1030 , \U1/keyexpantion/SB0/n752 ,
         \U1/keyexpantion/SB0/n707 , \U1/keyexpantion/SB0/n385 ;
  wire   [127:0] \U1/key ;
  wire   [7:0] \U1/rcon ;
  wire   [127:0] \U1/rkey ;
  wire   [127:0] \U1/rkey_next ;
  wire   [127:0] \U1/dat_next ;
  wire   [9:0] \U1/rnd ;
  wire   [31:0] \U1/aes_core/sc3 ;
  wire   [31:0] \U1/aes_core/sc2 ;
  wire   [31:0] \U1/aes_core/sc1 ;
  wire   [31:0] \U1/aes_core/sc0 ;
  wire   [31:0] \U1/aes_core/sb3 ;
  wire   [31:0] \U1/aes_core/sb2 ;
  wire   [31:0] \U1/aes_core/sb1 ;
  wire   [31:0] \U1/aes_core/sb0 ;
  wire   [31:0] \U1/keyexpantion/ws ;

  DFFNRPQ_X1M_A12TL trigger_reg ( .D(Dvld), .CKN(CLK), .R(N0), .Q(trigger) );
  DFFRPQ_X0P5M_A12TL KDrdy2_reg ( .D(Kvld), .CK(CLK), .R(N0), .Q(KDrdy2) );
  INV_X1M_A12TL U4 ( .A(RSTn), .Y(N0) );
  BUFH_X1M_A12TL \U1/U1103  ( .A(\U1/n1 ), .Y(\U1/n1108 ) );
  INV_X1M_A12TL \U1/U1102  ( .A(\U1/n1108 ), .Y(\U1/n1105 ) );
  INV_X1M_A12TL \U1/U1101  ( .A(\U1/n1108 ), .Y(\U1/n1104 ) );
  INV_X1M_A12TL \U1/U1100  ( .A(\U1/n1108 ), .Y(\U1/n1107 ) );
  INV_X1M_A12TL \U1/U1099  ( .A(\U1/n1108 ), .Y(\U1/n1106 ) );
  BUFH_X1M_A12TL \U1/U1098  ( .A(\U1/n1101 ), .Y(\U1/n1100 ) );
  BUFH_X1M_A12TL \U1/U1097  ( .A(\U1/n400 ), .Y(\U1/n1098 ) );
  BUFH_X1M_A12TL \U1/U1096  ( .A(\U1/n1097 ), .Y(\U1/n1095 ) );
  BUFH_X1M_A12TL \U1/U1095  ( .A(\U1/n1097 ), .Y(\U1/n1096 ) );
  BUFH_X1M_A12TL \U1/U1094  ( .A(\U1/n404 ), .Y(\U1/n670 ) );
  BUFH_X1M_A12TL \U1/U1093  ( .A(\U1/n5 ), .Y(\U1/n1103 ) );
  BUFH_X1M_A12TL \U1/U1092  ( .A(\U1/n7 ), .Y(\U1/n1099 ) );
  BUFH_X1M_A12TL \U1/U1091  ( .A(\U1/n5 ), .Y(\U1/n1102 ) );
  BUFH_X1M_A12TL \U1/U1090  ( .A(\U1/n6 ), .Y(\U1/n1101 ) );
  BUFH_X1M_A12TL \U1/U1089  ( .A(\U1/n402 ), .Y(\U1/n1097 ) );
  INV_X7P5M_A12TL \U1/U1073  ( .A(RSTn), .Y(\U1/rst ) );
  AND2_X1M_A12TL \U1/U1072  ( .A(KDrdy), .B(EN), .Y(\U1/n1 ) );
  INV_X1M_A12TL \U1/U922  ( .A(EN), .Y(\U1/n7 ) );
  NOR2_X1A_A12TL \U1/U3  ( .A(\U1/n1098 ), .B(KDrdy2), .Y(\U1/n404 ) );
  DFFRPQ_X2M_A12TL \U1/sel_reg  ( .D(\U1/n811 ), .CK(CLK), .R(\U1/rst ), .Q(
        \U1/sel ) );
  DFFRPQ_X0P5M_A12TL \U1/rnd_reg[9]  ( .D(\U1/n1085 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rnd [9]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[0]  ( .D(\U1/n948 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[0]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[1]  ( .D(\U1/n947 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[1]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[2]  ( .D(\U1/n946 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[2]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[3]  ( .D(\U1/n945 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[3]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[4]  ( .D(\U1/n944 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[4]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[5]  ( .D(\U1/n943 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[5]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[6]  ( .D(\U1/n942 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[6]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[7]  ( .D(\U1/n941 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[7]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[8]  ( .D(\U1/n940 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[8]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[9]  ( .D(\U1/n939 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[9]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[10]  ( .D(\U1/n938 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[10]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[11]  ( .D(\U1/n937 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[11]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[12]  ( .D(\U1/n936 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[12]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[13]  ( .D(\U1/n935 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[13]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[14]  ( .D(\U1/n934 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[14]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[15]  ( .D(\U1/n933 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[15]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[16]  ( .D(\U1/n932 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[16]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[17]  ( .D(\U1/n931 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[17]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[18]  ( .D(\U1/n930 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[18]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[19]  ( .D(\U1/n929 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[19]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[20]  ( .D(\U1/n928 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[20]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[21]  ( .D(\U1/n927 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[21]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[22]  ( .D(\U1/n926 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[22]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[23]  ( .D(\U1/n925 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[23]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[24]  ( .D(\U1/n924 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[24]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[25]  ( .D(\U1/n923 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[25]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[26]  ( .D(\U1/n922 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[26]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[27]  ( .D(\U1/n921 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[27]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[28]  ( .D(\U1/n920 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[28]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[29]  ( .D(\U1/n919 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[29]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[30]  ( .D(\U1/n918 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[30]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[31]  ( .D(\U1/n917 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[31]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[32]  ( .D(\U1/n916 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[32]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[33]  ( .D(\U1/n915 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[33]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[34]  ( .D(\U1/n914 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[34]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[35]  ( .D(\U1/n913 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[35]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[36]  ( .D(\U1/n912 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[36]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[37]  ( .D(\U1/n911 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[37]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[38]  ( .D(\U1/n910 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[38]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[39]  ( .D(\U1/n909 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[39]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[40]  ( .D(\U1/n908 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[40]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[41]  ( .D(\U1/n907 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[41]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[42]  ( .D(\U1/n906 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[42]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[43]  ( .D(\U1/n905 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[43]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[44]  ( .D(\U1/n904 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[44]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[45]  ( .D(\U1/n903 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[45]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[46]  ( .D(\U1/n902 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[46]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[47]  ( .D(\U1/n901 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[47]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[48]  ( .D(\U1/n900 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[48]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[49]  ( .D(\U1/n899 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[49]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[50]  ( .D(\U1/n898 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[50]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[51]  ( .D(\U1/n897 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[51]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[52]  ( .D(\U1/n896 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[52]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[53]  ( .D(\U1/n895 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[53]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[54]  ( .D(\U1/n894 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[54]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[55]  ( .D(\U1/n893 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[55]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[56]  ( .D(\U1/n892 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[56]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[57]  ( .D(\U1/n891 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[57]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[58]  ( .D(\U1/n890 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[58]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[59]  ( .D(\U1/n889 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[59]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[60]  ( .D(\U1/n888 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[60]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[61]  ( .D(\U1/n887 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[61]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[62]  ( .D(\U1/n886 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[62]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[63]  ( .D(\U1/n885 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[63]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[64]  ( .D(\U1/n884 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[64]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[65]  ( .D(\U1/n883 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[65]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[66]  ( .D(\U1/n882 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[66]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[67]  ( .D(\U1/n881 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[67]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[68]  ( .D(\U1/n880 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[68]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[69]  ( .D(\U1/n879 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[69]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[70]  ( .D(\U1/n878 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[70]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[71]  ( .D(\U1/n877 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[71]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[72]  ( .D(\U1/n876 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[72]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[73]  ( .D(\U1/n875 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[73]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[74]  ( .D(\U1/n874 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[74]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[75]  ( .D(\U1/n873 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[75]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[76]  ( .D(\U1/n872 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[76]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[77]  ( .D(\U1/n871 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[77]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[78]  ( .D(\U1/n870 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[78]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[79]  ( .D(\U1/n869 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[79]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[80]  ( .D(\U1/n868 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[80]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[81]  ( .D(\U1/n867 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[81]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[82]  ( .D(\U1/n866 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[82]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[83]  ( .D(\U1/n865 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[83]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[84]  ( .D(\U1/n864 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[84]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[85]  ( .D(\U1/n863 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[85]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[86]  ( .D(\U1/n862 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[86]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[87]  ( .D(\U1/n861 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[87]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[88]  ( .D(\U1/n860 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[88]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[89]  ( .D(\U1/n859 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[89]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[90]  ( .D(\U1/n858 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[90]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[91]  ( .D(\U1/n857 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[91]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[92]  ( .D(\U1/n856 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[92]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[93]  ( .D(\U1/n855 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[93]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[94]  ( .D(\U1/n854 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[94]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[95]  ( .D(\U1/n853 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[95]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[96]  ( .D(\U1/n852 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[96]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[97]  ( .D(\U1/n851 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[97]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[98]  ( .D(\U1/n850 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[98]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[99]  ( .D(\U1/n849 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[99]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[100]  ( .D(\U1/n848 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[100]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[101]  ( .D(\U1/n847 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[101]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[102]  ( .D(\U1/n846 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[102]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[103]  ( .D(\U1/n845 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[103]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[104]  ( .D(\U1/n844 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[104]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[105]  ( .D(\U1/n843 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[105]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[106]  ( .D(\U1/n842 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[106]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[107]  ( .D(\U1/n841 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[107]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[108]  ( .D(\U1/n840 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[108]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[109]  ( .D(\U1/n839 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[109]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[110]  ( .D(\U1/n838 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[110]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[111]  ( .D(\U1/n837 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[111]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[112]  ( .D(\U1/n836 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[112]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[113]  ( .D(\U1/n835 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[113]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[114]  ( .D(\U1/n834 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[114]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[115]  ( .D(\U1/n833 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[115]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[116]  ( .D(\U1/n832 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[116]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[64]  ( .D(\U1/n737 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [64]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[65]  ( .D(\U1/n736 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [65]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[66]  ( .D(\U1/n735 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [66]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[67]  ( .D(\U1/n734 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [67]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[68]  ( .D(\U1/n733 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [68]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[69]  ( .D(\U1/n732 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [69]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[70]  ( .D(\U1/n731 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [70]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[71]  ( .D(\U1/n730 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [71]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[72]  ( .D(\U1/n729 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [72]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[73]  ( .D(\U1/n728 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [73]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[74]  ( .D(\U1/n727 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [74]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[75]  ( .D(\U1/n726 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [75]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[76]  ( .D(\U1/n725 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [76]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[77]  ( .D(\U1/n724 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [77]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[32]  ( .D(\U1/n769 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [32]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[33]  ( .D(\U1/n768 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [33]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[34]  ( .D(\U1/n767 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [34]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[35]  ( .D(\U1/n766 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [35]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[36]  ( .D(\U1/n765 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [36]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[37]  ( .D(\U1/n764 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [37]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[38]  ( .D(\U1/n763 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [38]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[39]  ( .D(\U1/n762 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [39]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[40]  ( .D(\U1/n761 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [40]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[41]  ( .D(\U1/n760 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [41]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[42]  ( .D(\U1/n759 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [42]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[43]  ( .D(\U1/n758 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [43]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[44]  ( .D(\U1/n757 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [44]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[45]  ( .D(\U1/n756 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [45]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[46]  ( .D(\U1/n755 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [46]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[47]  ( .D(\U1/n754 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [47]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[48]  ( .D(\U1/n753 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [48]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[49]  ( .D(\U1/n752 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [49]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[50]  ( .D(\U1/n751 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [50]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[51]  ( .D(\U1/n750 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [51]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[52]  ( .D(\U1/n749 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [52]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[53]  ( .D(\U1/n748 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [53]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[54]  ( .D(\U1/n747 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [54]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[55]  ( .D(\U1/n746 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [55]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[56]  ( .D(\U1/n745 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [56]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[57]  ( .D(\U1/n744 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [57]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[58]  ( .D(\U1/n743 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [58]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[59]  ( .D(\U1/n742 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [59]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[60]  ( .D(\U1/n741 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [60]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[61]  ( .D(\U1/n740 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [61]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[62]  ( .D(\U1/n739 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [62]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[63]  ( .D(\U1/n738 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [63]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[6]  ( .D(\U1/n795 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [6]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[7]  ( .D(\U1/n794 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [7]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[8]  ( .D(\U1/n793 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [8]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[9]  ( .D(\U1/n792 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [9]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[10]  ( .D(\U1/n791 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [10]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[11]  ( .D(\U1/n790 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [11]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[12]  ( .D(\U1/n789 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [12]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[13]  ( .D(\U1/n788 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [13]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[14]  ( .D(\U1/n787 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [14]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[15]  ( .D(\U1/n786 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [15]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[16]  ( .D(\U1/n785 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [16]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[17]  ( .D(\U1/n784 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [17]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[18]  ( .D(\U1/n783 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [18]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[19]  ( .D(\U1/n782 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [19]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[20]  ( .D(\U1/n781 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [20]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[21]  ( .D(\U1/n780 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [21]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[22]  ( .D(\U1/n779 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [22]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[23]  ( .D(\U1/n778 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [23]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[24]  ( .D(\U1/n777 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [24]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[25]  ( .D(\U1/n776 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [25]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[26]  ( .D(\U1/n775 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [26]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[27]  ( .D(\U1/n774 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [27]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[28]  ( .D(\U1/n773 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [28]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[29]  ( .D(\U1/n772 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [29]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[30]  ( .D(\U1/n771 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [30]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[31]  ( .D(\U1/n770 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [31]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[0]  ( .D(\U1/n801 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [0]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[1]  ( .D(\U1/n800 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [1]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[2]  ( .D(\U1/n799 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [2]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[3]  ( .D(\U1/n798 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [3]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[4]  ( .D(\U1/n797 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [4]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[5]  ( .D(\U1/n796 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [5]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[78]  ( .D(\U1/n723 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [78]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[79]  ( .D(\U1/n722 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [79]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[80]  ( .D(\U1/n721 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [80]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[81]  ( .D(\U1/n720 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [81]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[82]  ( .D(\U1/n719 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [82]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[83]  ( .D(\U1/n718 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [83]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[84]  ( .D(\U1/n717 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [84]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[85]  ( .D(\U1/n716 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [85]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[86]  ( .D(\U1/n715 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [86]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[87]  ( .D(\U1/n714 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [87]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[88]  ( .D(\U1/n713 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [88]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[89]  ( .D(\U1/n712 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [89]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[90]  ( .D(\U1/n711 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [90]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[91]  ( .D(\U1/n710 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [91]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[92]  ( .D(\U1/n709 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [92]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[93]  ( .D(\U1/n708 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [93]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[94]  ( .D(\U1/n707 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [94]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[95]  ( .D(\U1/n706 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [95]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[96]  ( .D(\U1/n705 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [96]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[97]  ( .D(\U1/n704 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [97]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[98]  ( .D(\U1/n703 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [98]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[99]  ( .D(\U1/n702 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rkey [99]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[100]  ( .D(\U1/n701 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [100]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[101]  ( .D(\U1/n700 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [101]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[102]  ( .D(\U1/n699 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [102]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[103]  ( .D(\U1/n698 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [103]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[104]  ( .D(\U1/n697 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [104]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[105]  ( .D(\U1/n696 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [105]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[106]  ( .D(\U1/n695 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [106]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[107]  ( .D(\U1/n694 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [107]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[108]  ( .D(\U1/n693 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [108]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[109]  ( .D(\U1/n692 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [109]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[110]  ( .D(\U1/n691 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [110]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[111]  ( .D(\U1/n690 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [111]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[112]  ( .D(\U1/n689 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [112]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[113]  ( .D(\U1/n688 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [113]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[114]  ( .D(\U1/n687 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [114]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[115]  ( .D(\U1/n686 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [115]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[116]  ( .D(\U1/n685 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [116]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[117]  ( .D(\U1/n831 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[117]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[118]  ( .D(\U1/n830 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[118]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[119]  ( .D(\U1/n829 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[119]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[120]  ( .D(\U1/n828 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[120]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[121]  ( .D(\U1/n827 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[121]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[122]  ( .D(\U1/n826 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[122]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[123]  ( .D(\U1/n825 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[123]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[124]  ( .D(\U1/n824 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[124]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[125]  ( .D(\U1/n823 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[125]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[126]  ( .D(\U1/n822 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[126]) );
  DFFRPQ_X0P5M_A12TL \U1/dat_reg[127]  ( .D(\U1/n821 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dout[127]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[117]  ( .D(\U1/n684 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [117]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[118]  ( .D(\U1/n683 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [118]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[119]  ( .D(\U1/n682 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [119]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[120]  ( .D(\U1/n681 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [120]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[121]  ( .D(\U1/n680 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [121]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[127]  ( .D(\U1/n674 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [127]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[122]  ( .D(\U1/n679 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [122]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[123]  ( .D(\U1/n678 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [123]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[124]  ( .D(\U1/n677 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [124]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[125]  ( .D(\U1/n676 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [125]) );
  DFFRPQ_X0P5M_A12TL \U1/rkey_reg[126]  ( .D(\U1/n675 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/rkey [126]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[44]  ( .D(\U1/n1001 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [44]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[45]  ( .D(\U1/n1002 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [45]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[46]  ( .D(\U1/n1003 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [46]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[47]  ( .D(\U1/n1004 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [47]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[48]  ( .D(\U1/n1005 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [48]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[49]  ( .D(\U1/n1006 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [49]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[50]  ( .D(\U1/n1007 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [50]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[51]  ( .D(\U1/n1008 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [51]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[52]  ( .D(\U1/n1009 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [52]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[53]  ( .D(\U1/n1010 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [53]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[54]  ( .D(\U1/n1011 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [54]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[55]  ( .D(\U1/n1012 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [55]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[56]  ( .D(\U1/n1013 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [56]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[57]  ( .D(\U1/n1014 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [57]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[58]  ( .D(\U1/n1015 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [58]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[59]  ( .D(\U1/n1016 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [59]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[60]  ( .D(\U1/n1017 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [60]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[61]  ( .D(\U1/n1018 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [61]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[62]  ( .D(\U1/n1019 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [62]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[63]  ( .D(\U1/n1020 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [63]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[64]  ( .D(\U1/n1021 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [64]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[65]  ( .D(\U1/n1022 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [65]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[66]  ( .D(\U1/n1023 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [66]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[67]  ( .D(\U1/n1024 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [67]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[68]  ( .D(\U1/n1025 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [68]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[69]  ( .D(\U1/n1026 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [69]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[70]  ( .D(\U1/n1027 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [70]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[71]  ( .D(\U1/n1028 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [71]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[72]  ( .D(\U1/n1029 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [72]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[73]  ( .D(\U1/n1030 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [73]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[74]  ( .D(\U1/n1031 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [74]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[75]  ( .D(\U1/n1032 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [75]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[76]  ( .D(\U1/n1033 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [76]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[77]  ( .D(\U1/n1034 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [77]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[78]  ( .D(\U1/n1035 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [78]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[79]  ( .D(\U1/n1036 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [79]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[80]  ( .D(\U1/n1037 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [80]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[81]  ( .D(\U1/n1038 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [81]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[82]  ( .D(\U1/n1039 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [82]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[83]  ( .D(\U1/n1040 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [83]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[84]  ( .D(\U1/n1041 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [84]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[85]  ( .D(\U1/n1042 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [85]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[86]  ( .D(\U1/n1043 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [86]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[87]  ( .D(\U1/n1044 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [87]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[88]  ( .D(\U1/n1045 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [88]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[89]  ( .D(\U1/n1046 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [89]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[90]  ( .D(\U1/n1047 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [90]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[91]  ( .D(\U1/n1048 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [91]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[92]  ( .D(\U1/n1049 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [92]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[93]  ( .D(\U1/n1050 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [93]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[94]  ( .D(\U1/n1051 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [94]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[95]  ( .D(\U1/n1052 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [95]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[96]  ( .D(\U1/n1053 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [96]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[97]  ( .D(\U1/n1054 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [97]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[98]  ( .D(\U1/n1055 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [98]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[99]  ( .D(\U1/n1056 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [99]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[100]  ( .D(\U1/n1057 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [100]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[101]  ( .D(\U1/n1058 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [101]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[102]  ( .D(\U1/n1059 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [102]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[103]  ( .D(\U1/n1060 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [103]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[104]  ( .D(\U1/n1061 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [104]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[105]  ( .D(\U1/n1062 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [105]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[106]  ( .D(\U1/n1063 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [106]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[0]  ( .D(\U1/n957 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [0]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[1]  ( .D(\U1/n958 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [1]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[2]  ( .D(\U1/n959 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [2]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[3]  ( .D(\U1/n960 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [3]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[4]  ( .D(\U1/n961 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [4]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[5]  ( .D(\U1/n962 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [5]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[6]  ( .D(\U1/n963 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [6]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[7]  ( .D(\U1/n964 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [7]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[8]  ( .D(\U1/n965 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [8]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[9]  ( .D(\U1/n966 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [9]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[10]  ( .D(\U1/n967 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [10]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[11]  ( .D(\U1/n968 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [11]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[12]  ( .D(\U1/n969 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [12]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[13]  ( .D(\U1/n970 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [13]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[14]  ( .D(\U1/n971 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [14]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[15]  ( .D(\U1/n972 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [15]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[16]  ( .D(\U1/n973 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [16]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[17]  ( .D(\U1/n974 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [17]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[18]  ( .D(\U1/n975 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [18]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[19]  ( .D(\U1/n976 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [19]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[20]  ( .D(\U1/n977 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [20]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[21]  ( .D(\U1/n978 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [21]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[22]  ( .D(\U1/n979 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [22]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[23]  ( .D(\U1/n980 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [23]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[24]  ( .D(\U1/n981 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [24]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[25]  ( .D(\U1/n982 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [25]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[26]  ( .D(\U1/n983 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [26]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[27]  ( .D(\U1/n984 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [27]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[28]  ( .D(\U1/n985 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [28]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[29]  ( .D(\U1/n986 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [29]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[30]  ( .D(\U1/n987 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [30]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[31]  ( .D(\U1/n988 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [31]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[32]  ( .D(\U1/n989 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [32]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[33]  ( .D(\U1/n990 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [33]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[34]  ( .D(\U1/n991 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [34]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[35]  ( .D(\U1/n992 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [35]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[36]  ( .D(\U1/n993 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [36]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[37]  ( .D(\U1/n994 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [37]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[38]  ( .D(\U1/n995 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [38]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[39]  ( .D(\U1/n996 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [39]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[40]  ( .D(\U1/n997 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [40]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[41]  ( .D(\U1/n998 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [41]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[42]  ( .D(\U1/n999 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [42]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[43]  ( .D(\U1/n1000 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/key [43]) );
  DFFRPQ_X0P5M_A12TL \U1/rcon_reg[7]  ( .D(\U1/n949 ), .CK(CLK), .R(\U1/rst ), 
        .Q(\U1/rcon [7]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[107]  ( .D(\U1/n1064 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [107]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[108]  ( .D(\U1/n1065 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [108]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[109]  ( .D(\U1/n1066 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [109]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[110]  ( .D(\U1/n1067 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [110]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[111]  ( .D(\U1/n1068 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [111]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[112]  ( .D(\U1/n1069 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [112]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[113]  ( .D(\U1/n1070 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [113]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[114]  ( .D(\U1/n1071 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [114]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[115]  ( .D(\U1/n1072 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [115]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[116]  ( .D(\U1/n1073 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [116]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[117]  ( .D(\U1/n1074 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [117]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[118]  ( .D(\U1/n1075 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [118]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[127]  ( .D(\U1/n1084 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [127]) );
  DFFRPQ_X0P5M_A12TL \U1/BSY_reg  ( .D(\U1/n809 ), .CK(CLK), .R(\U1/rst ), .Q(
        BSY) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[119]  ( .D(\U1/n1076 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [119]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[120]  ( .D(\U1/n1077 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [120]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[121]  ( .D(\U1/n1078 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [121]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[122]  ( .D(\U1/n1079 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [122]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[123]  ( .D(\U1/n1080 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [123]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[124]  ( .D(\U1/n1081 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [124]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[125]  ( .D(\U1/n1082 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [125]) );
  DFFRPQ_X0P5M_A12TL \U1/key_reg[126]  ( .D(\U1/n1083 ), .CK(CLK), .R(\U1/rst ), .Q(\U1/key [126]) );
  DFFRPQ_X0P5M_A12TL \U1/Kvld_reg  ( .D(\U1/n820 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Kvld) );
  DFFRPQ_X0P5M_A12TL \U1/Dvld_reg  ( .D(\U1/n810 ), .CK(CLK), .R(\U1/rst ), 
        .Q(Dvld) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[2]  ( .D(\U1/n1092 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n818 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[3]  ( .D(\U1/n1091 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n817 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[4]  ( .D(\U1/n1090 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n816 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[5]  ( .D(\U1/n1089 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n815 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[6]  ( .D(\U1/n1088 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n814 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[7]  ( .D(\U1/n1087 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n813 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[8]  ( .D(\U1/n1086 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n812 ) );
  DFFRPQN_X1M_A12TL \U1/rnd_reg[1]  ( .D(\U1/n1093 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n819 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[2]  ( .D(\U1/n954 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n806 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[5]  ( .D(\U1/n951 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n803 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[6]  ( .D(\U1/n950 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n802 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[1]  ( .D(\U1/n955 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n807 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[3]  ( .D(\U1/n953 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n805 ) );
  DFFRPQN_X1M_A12TL \U1/rcon_reg[4]  ( .D(\U1/n952 ), .CK(CLK), .R(\U1/rst ), 
        .QN(\U1/n804 ) );
  DFFSQN_X1M_A12TL \U1/rcon_reg[0]  ( .D(\U1/n956 ), .CK(CLK), .SN(RSTn), .QN(
        \U1/n808 ) );
  DFFSQ_X1M_A12TL \U1/rnd_reg[0]  ( .D(\U1/n1094 ), .CK(CLK), .SN(RSTn), .Q(
        \U1/rnd [0]) );
  NAND2_X0P5A_A12TL \U1/U1088  ( .A(KDrdy2), .B(EN), .Y(\U1/n661 ) );
  OAI21_X0P5M_A12TL \U1/U1087  ( .A0(\U1/rnd [0]), .A1(\U1/n1099 ), .B0(
        \U1/n661 ), .Y(\U1/n673 ) );
  INV_X0P5B_A12TL \U1/U1086  ( .A(\U1/n673 ), .Y(\U1/n671 ) );
  INV_X0P5B_A12TL \U1/U1085  ( .A(\U1/rnd [9]), .Y(\U1/n672 ) );
  INV_X0P5B_A12TL \U1/U1084  ( .A(\U1/rnd [0]), .Y(\U1/n389 ) );
  OAI22_X0P5M_A12TL \U1/U1083  ( .A0(\U1/n671 ), .A1(\U1/n672 ), .B0(\U1/n389 ), .B1(\U1/n673 ), .Y(\U1/n1094 ) );
  OAI22_X0P5M_A12TL \U1/U1082  ( .A0(\U1/n671 ), .A1(\U1/n389 ), .B0(\U1/n819 ), .B1(\U1/n673 ), .Y(\U1/n1093 ) );
  OAI22_X0P5M_A12TL \U1/U1081  ( .A0(\U1/n819 ), .A1(\U1/n671 ), .B0(\U1/n818 ), .B1(\U1/n673 ), .Y(\U1/n1092 ) );
  OAI22_X0P5M_A12TL \U1/U1080  ( .A0(\U1/n818 ), .A1(\U1/n671 ), .B0(\U1/n817 ), .B1(\U1/n673 ), .Y(\U1/n1091 ) );
  OAI22_X0P5M_A12TL \U1/U1079  ( .A0(\U1/n817 ), .A1(\U1/n671 ), .B0(\U1/n816 ), .B1(\U1/n673 ), .Y(\U1/n1090 ) );
  OAI22_X0P5M_A12TL \U1/U1078  ( .A0(\U1/n816 ), .A1(\U1/n671 ), .B0(\U1/n815 ), .B1(\U1/n673 ), .Y(\U1/n1089 ) );
  OAI22_X0P5M_A12TL \U1/U1077  ( .A0(\U1/n815 ), .A1(\U1/n671 ), .B0(\U1/n814 ), .B1(\U1/n673 ), .Y(\U1/n1088 ) );
  OAI22_X0P5M_A12TL \U1/U1076  ( .A0(\U1/n814 ), .A1(\U1/n671 ), .B0(\U1/n813 ), .B1(\U1/n673 ), .Y(\U1/n1087 ) );
  OAI22_X0P5M_A12TL \U1/U1075  ( .A0(\U1/n813 ), .A1(\U1/n671 ), .B0(\U1/n812 ), .B1(\U1/n673 ), .Y(\U1/n1086 ) );
  OAI22_X0P5M_A12TL \U1/U1074  ( .A0(\U1/n812 ), .A1(\U1/n671 ), .B0(\U1/n672 ), .B1(\U1/n673 ), .Y(\U1/n1085 ) );
  AO22_X0P5M_A12TL \U1/U1071  ( .A0(\U1/n1104 ), .A1(\U1/key [127]), .B0(
        \U1/n1108 ), .B1(Kin[127]), .Y(\U1/n1084 ) );
  AO22_X0P5M_A12TL \U1/U1070  ( .A0(\U1/n1104 ), .A1(\U1/key [126]), .B0(
        \U1/n1108 ), .B1(Kin[126]), .Y(\U1/n1083 ) );
  AO22_X0P5M_A12TL \U1/U1069  ( .A0(\U1/n1105 ), .A1(\U1/key [125]), .B0(
        \U1/n1108 ), .B1(Kin[125]), .Y(\U1/n1082 ) );
  AO22_X0P5M_A12TL \U1/U1068  ( .A0(\U1/n1106 ), .A1(\U1/key [124]), .B0(
        \U1/n1108 ), .B1(Kin[124]), .Y(\U1/n1081 ) );
  AO22_X0P5M_A12TL \U1/U1067  ( .A0(\U1/n1106 ), .A1(\U1/key [123]), .B0(
        \U1/n1108 ), .B1(Kin[123]), .Y(\U1/n1080 ) );
  AO22_X0P5M_A12TL \U1/U1066  ( .A0(\U1/n1104 ), .A1(\U1/key [122]), .B0(
        \U1/n1108 ), .B1(Kin[122]), .Y(\U1/n1079 ) );
  AO22_X0P5M_A12TL \U1/U1065  ( .A0(\U1/n1107 ), .A1(\U1/key [121]), .B0(
        \U1/n1108 ), .B1(Kin[121]), .Y(\U1/n1078 ) );
  AO22_X0P5M_A12TL \U1/U1064  ( .A0(\U1/n1104 ), .A1(\U1/key [120]), .B0(
        \U1/n1108 ), .B1(Kin[120]), .Y(\U1/n1077 ) );
  AO22_X0P5M_A12TL \U1/U1063  ( .A0(\U1/n1105 ), .A1(\U1/key [119]), .B0(
        \U1/n1108 ), .B1(Kin[119]), .Y(\U1/n1076 ) );
  AO22_X0P5M_A12TL \U1/U1062  ( .A0(\U1/n1107 ), .A1(\U1/key [118]), .B0(
        \U1/n1108 ), .B1(Kin[118]), .Y(\U1/n1075 ) );
  AO22_X0P5M_A12TL \U1/U1061  ( .A0(\U1/n1106 ), .A1(\U1/key [117]), .B0(
        \U1/n1108 ), .B1(Kin[117]), .Y(\U1/n1074 ) );
  AO22_X0P5M_A12TL \U1/U1060  ( .A0(\U1/n1106 ), .A1(\U1/key [116]), .B0(
        \U1/n1108 ), .B1(Kin[116]), .Y(\U1/n1073 ) );
  AO22_X0P5M_A12TL \U1/U1059  ( .A0(\U1/n1104 ), .A1(\U1/key [115]), .B0(
        \U1/n1108 ), .B1(Kin[115]), .Y(\U1/n1072 ) );
  AO22_X0P5M_A12TL \U1/U1058  ( .A0(\U1/n1107 ), .A1(\U1/key [114]), .B0(
        \U1/n1108 ), .B1(Kin[114]), .Y(\U1/n1071 ) );
  AO22_X0P5M_A12TL \U1/U1057  ( .A0(\U1/n1104 ), .A1(\U1/key [113]), .B0(
        \U1/n1108 ), .B1(Kin[113]), .Y(\U1/n1070 ) );
  AO22_X0P5M_A12TL \U1/U1056  ( .A0(\U1/n1106 ), .A1(\U1/key [112]), .B0(
        \U1/n1108 ), .B1(Kin[112]), .Y(\U1/n1069 ) );
  AO22_X0P5M_A12TL \U1/U1055  ( .A0(\U1/n1105 ), .A1(\U1/key [111]), .B0(
        \U1/n1108 ), .B1(Kin[111]), .Y(\U1/n1068 ) );
  AO22_X0P5M_A12TL \U1/U1054  ( .A0(\U1/n1106 ), .A1(\U1/key [110]), .B0(
        \U1/n1108 ), .B1(Kin[110]), .Y(\U1/n1067 ) );
  AO22_X0P5M_A12TL \U1/U1053  ( .A0(\U1/n1104 ), .A1(\U1/key [109]), .B0(
        \U1/n1108 ), .B1(Kin[109]), .Y(\U1/n1066 ) );
  AO22_X0P5M_A12TL \U1/U1052  ( .A0(\U1/n1105 ), .A1(\U1/key [108]), .B0(
        \U1/n1108 ), .B1(Kin[108]), .Y(\U1/n1065 ) );
  AO22_X0P5M_A12TL \U1/U1051  ( .A0(\U1/n1105 ), .A1(\U1/key [107]), .B0(
        \U1/n1108 ), .B1(Kin[107]), .Y(\U1/n1064 ) );
  AO22_X0P5M_A12TL \U1/U1050  ( .A0(\U1/n1107 ), .A1(\U1/key [106]), .B0(
        \U1/n1108 ), .B1(Kin[106]), .Y(\U1/n1063 ) );
  AO22_X0P5M_A12TL \U1/U1049  ( .A0(\U1/n1106 ), .A1(\U1/key [105]), .B0(
        \U1/n1 ), .B1(Kin[105]), .Y(\U1/n1062 ) );
  AO22_X0P5M_A12TL \U1/U1048  ( .A0(\U1/n1106 ), .A1(\U1/key [104]), .B0(
        \U1/n1 ), .B1(Kin[104]), .Y(\U1/n1061 ) );
  AO22_X0P5M_A12TL \U1/U1047  ( .A0(\U1/n1104 ), .A1(\U1/key [103]), .B0(
        \U1/n1108 ), .B1(Kin[103]), .Y(\U1/n1060 ) );
  AO22_X0P5M_A12TL \U1/U1046  ( .A0(\U1/n1107 ), .A1(\U1/key [102]), .B0(
        \U1/n1 ), .B1(Kin[102]), .Y(\U1/n1059 ) );
  AO22_X0P5M_A12TL \U1/U1045  ( .A0(\U1/n1106 ), .A1(\U1/key [101]), .B0(
        \U1/n1108 ), .B1(Kin[101]), .Y(\U1/n1058 ) );
  AO22_X0P5M_A12TL \U1/U1044  ( .A0(\U1/n1107 ), .A1(\U1/key [100]), .B0(
        \U1/n1108 ), .B1(Kin[100]), .Y(\U1/n1057 ) );
  AO22_X0P5M_A12TL \U1/U1043  ( .A0(\U1/n1105 ), .A1(\U1/key [99]), .B0(
        \U1/n1108 ), .B1(Kin[99]), .Y(\U1/n1056 ) );
  AO22_X0P5M_A12TL \U1/U1042  ( .A0(\U1/n1107 ), .A1(\U1/key [98]), .B0(
        \U1/n1108 ), .B1(Kin[98]), .Y(\U1/n1055 ) );
  AO22_X0P5M_A12TL \U1/U1041  ( .A0(\U1/n1107 ), .A1(\U1/key [97]), .B0(
        \U1/n1108 ), .B1(Kin[97]), .Y(\U1/n1054 ) );
  AO22_X0P5M_A12TL \U1/U1040  ( .A0(\U1/n1106 ), .A1(\U1/key [96]), .B0(
        \U1/n1108 ), .B1(Kin[96]), .Y(\U1/n1053 ) );
  AO22_X0P5M_A12TL \U1/U1039  ( .A0(\U1/n1106 ), .A1(\U1/key [95]), .B0(
        \U1/n1108 ), .B1(Kin[95]), .Y(\U1/n1052 ) );
  AO22_X0P5M_A12TL \U1/U1038  ( .A0(\U1/n1107 ), .A1(\U1/key [94]), .B0(
        \U1/n1 ), .B1(Kin[94]), .Y(\U1/n1051 ) );
  AO22_X0P5M_A12TL \U1/U1037  ( .A0(\U1/n1106 ), .A1(\U1/key [93]), .B0(
        \U1/n1 ), .B1(Kin[93]), .Y(\U1/n1050 ) );
  AO22_X0P5M_A12TL \U1/U1036  ( .A0(\U1/n1104 ), .A1(\U1/key [92]), .B0(
        \U1/n1 ), .B1(Kin[92]), .Y(\U1/n1049 ) );
  AO22_X0P5M_A12TL \U1/U1035  ( .A0(\U1/n1105 ), .A1(\U1/key [91]), .B0(
        \U1/n1 ), .B1(Kin[91]), .Y(\U1/n1048 ) );
  AO22_X0P5M_A12TL \U1/U1034  ( .A0(\U1/n1107 ), .A1(\U1/key [90]), .B0(
        \U1/n1 ), .B1(Kin[90]), .Y(\U1/n1047 ) );
  AO22_X0P5M_A12TL \U1/U1033  ( .A0(\U1/n1107 ), .A1(\U1/key [89]), .B0(
        \U1/n1 ), .B1(Kin[89]), .Y(\U1/n1046 ) );
  AO22_X0P5M_A12TL \U1/U1032  ( .A0(\U1/n1107 ), .A1(\U1/key [88]), .B0(
        \U1/n1108 ), .B1(Kin[88]), .Y(\U1/n1045 ) );
  AO22_X0P5M_A12TL \U1/U1031  ( .A0(\U1/n1105 ), .A1(\U1/key [87]), .B0(
        \U1/n1 ), .B1(Kin[87]), .Y(\U1/n1044 ) );
  AO22_X0P5M_A12TL \U1/U1030  ( .A0(\U1/n1107 ), .A1(\U1/key [86]), .B0(
        \U1/n1 ), .B1(Kin[86]), .Y(\U1/n1043 ) );
  AO22_X0P5M_A12TL \U1/U1029  ( .A0(\U1/n1106 ), .A1(\U1/key [85]), .B0(
        \U1/n1 ), .B1(Kin[85]), .Y(\U1/n1042 ) );
  AO22_X0P5M_A12TL \U1/U1028  ( .A0(\U1/n1106 ), .A1(\U1/key [84]), .B0(
        \U1/n1 ), .B1(Kin[84]), .Y(\U1/n1041 ) );
  AO22_X0P5M_A12TL \U1/U1027  ( .A0(\U1/n1104 ), .A1(\U1/key [83]), .B0(
        \U1/n1 ), .B1(Kin[83]), .Y(\U1/n1040 ) );
  AO22_X0P5M_A12TL \U1/U1026  ( .A0(\U1/n1104 ), .A1(\U1/key [82]), .B0(
        \U1/n1 ), .B1(Kin[82]), .Y(\U1/n1039 ) );
  AO22_X0P5M_A12TL \U1/U1025  ( .A0(\U1/n1104 ), .A1(\U1/key [81]), .B0(
        \U1/n1 ), .B1(Kin[81]), .Y(\U1/n1038 ) );
  AO22_X0P5M_A12TL \U1/U1024  ( .A0(\U1/n1106 ), .A1(\U1/key [80]), .B0(
        \U1/n1 ), .B1(Kin[80]), .Y(\U1/n1037 ) );
  AO22_X0P5M_A12TL \U1/U1023  ( .A0(\U1/n1105 ), .A1(\U1/key [79]), .B0(
        \U1/n1 ), .B1(Kin[79]), .Y(\U1/n1036 ) );
  AO22_X0P5M_A12TL \U1/U1022  ( .A0(\U1/n1106 ), .A1(\U1/key [78]), .B0(
        \U1/n1 ), .B1(Kin[78]), .Y(\U1/n1035 ) );
  AO22_X0P5M_A12TL \U1/U1021  ( .A0(\U1/n1107 ), .A1(\U1/key [77]), .B0(
        \U1/n1 ), .B1(Kin[77]), .Y(\U1/n1034 ) );
  AO22_X0P5M_A12TL \U1/U1020  ( .A0(\U1/n1107 ), .A1(\U1/key [76]), .B0(
        \U1/n1 ), .B1(Kin[76]), .Y(\U1/n1033 ) );
  AO22_X0P5M_A12TL \U1/U1019  ( .A0(\U1/n1104 ), .A1(\U1/key [75]), .B0(
        \U1/n1 ), .B1(Kin[75]), .Y(\U1/n1032 ) );
  AO22_X0P5M_A12TL \U1/U1018  ( .A0(\U1/n1105 ), .A1(\U1/key [74]), .B0(
        \U1/n1 ), .B1(Kin[74]), .Y(\U1/n1031 ) );
  AO22_X0P5M_A12TL \U1/U1017  ( .A0(\U1/n1104 ), .A1(\U1/key [73]), .B0(
        \U1/n1 ), .B1(Kin[73]), .Y(\U1/n1030 ) );
  AO22_X0P5M_A12TL \U1/U1016  ( .A0(\U1/n1107 ), .A1(\U1/key [72]), .B0(
        \U1/n1 ), .B1(Kin[72]), .Y(\U1/n1029 ) );
  AO22_X0P5M_A12TL \U1/U1015  ( .A0(\U1/n1105 ), .A1(\U1/key [71]), .B0(
        \U1/n1 ), .B1(Kin[71]), .Y(\U1/n1028 ) );
  AO22_X0P5M_A12TL \U1/U1014  ( .A0(\U1/n1106 ), .A1(\U1/key [70]), .B0(
        \U1/n1108 ), .B1(Kin[70]), .Y(\U1/n1027 ) );
  AO22_X0P5M_A12TL \U1/U1013  ( .A0(\U1/n1106 ), .A1(\U1/key [69]), .B0(
        \U1/n1 ), .B1(Kin[69]), .Y(\U1/n1026 ) );
  AO22_X0P5M_A12TL \U1/U1012  ( .A0(\U1/n1106 ), .A1(\U1/key [68]), .B0(
        \U1/n1 ), .B1(Kin[68]), .Y(\U1/n1025 ) );
  AO22_X0P5M_A12TL \U1/U1011  ( .A0(\U1/n1106 ), .A1(\U1/key [67]), .B0(
        \U1/n1 ), .B1(Kin[67]), .Y(\U1/n1024 ) );
  AO22_X0P5M_A12TL \U1/U1010  ( .A0(\U1/n1107 ), .A1(\U1/key [66]), .B0(
        \U1/n1 ), .B1(Kin[66]), .Y(\U1/n1023 ) );
  AO22_X0P5M_A12TL \U1/U1009  ( .A0(\U1/n1107 ), .A1(\U1/key [65]), .B0(
        \U1/n1 ), .B1(Kin[65]), .Y(\U1/n1022 ) );
  AO22_X0P5M_A12TL \U1/U1008  ( .A0(\U1/n1104 ), .A1(\U1/key [64]), .B0(
        \U1/n1 ), .B1(Kin[64]), .Y(\U1/n1021 ) );
  AO22_X0P5M_A12TL \U1/U1007  ( .A0(\U1/n1105 ), .A1(\U1/key [63]), .B0(
        \U1/n1 ), .B1(Kin[63]), .Y(\U1/n1020 ) );
  AO22_X0P5M_A12TL \U1/U1006  ( .A0(\U1/n1107 ), .A1(\U1/key [62]), .B0(
        \U1/n1 ), .B1(Kin[62]), .Y(\U1/n1019 ) );
  AO22_X0P5M_A12TL \U1/U1005  ( .A0(\U1/n1106 ), .A1(\U1/key [61]), .B0(
        \U1/n1 ), .B1(Kin[61]), .Y(\U1/n1018 ) );
  AO22_X0P5M_A12TL \U1/U1004  ( .A0(\U1/n1105 ), .A1(\U1/key [60]), .B0(
        \U1/n1 ), .B1(Kin[60]), .Y(\U1/n1017 ) );
  AO22_X0P5M_A12TL \U1/U1003  ( .A0(\U1/n1106 ), .A1(\U1/key [59]), .B0(
        \U1/n1 ), .B1(Kin[59]), .Y(\U1/n1016 ) );
  AO22_X0P5M_A12TL \U1/U1002  ( .A0(\U1/n1105 ), .A1(\U1/key [58]), .B0(
        \U1/n1 ), .B1(Kin[58]), .Y(\U1/n1015 ) );
  AO22_X0P5M_A12TL \U1/U1001  ( .A0(\U1/n1107 ), .A1(\U1/key [57]), .B0(
        \U1/n1 ), .B1(Kin[57]), .Y(\U1/n1014 ) );
  AO22_X0P5M_A12TL \U1/U1000  ( .A0(\U1/n1106 ), .A1(\U1/key [56]), .B0(
        \U1/n1 ), .B1(Kin[56]), .Y(\U1/n1013 ) );
  AO22_X0P5M_A12TL \U1/U999  ( .A0(\U1/n1104 ), .A1(\U1/key [55]), .B0(\U1/n1 ), .B1(Kin[55]), .Y(\U1/n1012 ) );
  AO22_X0P5M_A12TL \U1/U998  ( .A0(\U1/n1104 ), .A1(\U1/key [54]), .B0(\U1/n1 ), .B1(Kin[54]), .Y(\U1/n1011 ) );
  AO22_X0P5M_A12TL \U1/U997  ( .A0(\U1/n1105 ), .A1(\U1/key [53]), .B0(\U1/n1 ), .B1(Kin[53]), .Y(\U1/n1010 ) );
  AO22_X0P5M_A12TL \U1/U996  ( .A0(\U1/n1107 ), .A1(\U1/key [52]), .B0(
        \U1/n1108 ), .B1(Kin[52]), .Y(\U1/n1009 ) );
  AO22_X0P5M_A12TL \U1/U995  ( .A0(\U1/n1105 ), .A1(\U1/key [51]), .B0(\U1/n1 ), .B1(Kin[51]), .Y(\U1/n1008 ) );
  AO22_X0P5M_A12TL \U1/U994  ( .A0(\U1/n1107 ), .A1(\U1/key [50]), .B0(\U1/n1 ), .B1(Kin[50]), .Y(\U1/n1007 ) );
  AO22_X0P5M_A12TL \U1/U993  ( .A0(\U1/n1106 ), .A1(\U1/key [49]), .B0(\U1/n1 ), .B1(Kin[49]), .Y(\U1/n1006 ) );
  AO22_X0P5M_A12TL \U1/U992  ( .A0(\U1/n1104 ), .A1(\U1/key [48]), .B0(\U1/n1 ), .B1(Kin[48]), .Y(\U1/n1005 ) );
  AO22_X0P5M_A12TL \U1/U991  ( .A0(\U1/n1106 ), .A1(\U1/key [47]), .B0(\U1/n1 ), .B1(Kin[47]), .Y(\U1/n1004 ) );
  AO22_X0P5M_A12TL \U1/U990  ( .A0(\U1/n1105 ), .A1(\U1/key [46]), .B0(\U1/n1 ), .B1(Kin[46]), .Y(\U1/n1003 ) );
  AO22_X0P5M_A12TL \U1/U989  ( .A0(\U1/n1105 ), .A1(\U1/key [45]), .B0(\U1/n1 ), .B1(Kin[45]), .Y(\U1/n1002 ) );
  AO22_X0P5M_A12TL \U1/U988  ( .A0(\U1/n1104 ), .A1(\U1/key [44]), .B0(\U1/n1 ), .B1(Kin[44]), .Y(\U1/n1001 ) );
  AO22_X0P5M_A12TL \U1/U987  ( .A0(\U1/n1107 ), .A1(\U1/key [43]), .B0(\U1/n1 ), .B1(Kin[43]), .Y(\U1/n1000 ) );
  AO22_X0P5M_A12TL \U1/U986  ( .A0(\U1/n1104 ), .A1(\U1/key [42]), .B0(\U1/n1 ), .B1(Kin[42]), .Y(\U1/n999 ) );
  AO22_X0P5M_A12TL \U1/U985  ( .A0(\U1/n1107 ), .A1(\U1/key [41]), .B0(\U1/n1 ), .B1(Kin[41]), .Y(\U1/n998 ) );
  AO22_X0P5M_A12TL \U1/U984  ( .A0(\U1/n1106 ), .A1(\U1/key [40]), .B0(\U1/n1 ), .B1(Kin[40]), .Y(\U1/n997 ) );
  AO22_X0P5M_A12TL \U1/U983  ( .A0(\U1/n1105 ), .A1(\U1/key [39]), .B0(\U1/n1 ), .B1(Kin[39]), .Y(\U1/n996 ) );
  AO22_X0P5M_A12TL \U1/U982  ( .A0(\U1/n1106 ), .A1(\U1/key [38]), .B0(\U1/n1 ), .B1(Kin[38]), .Y(\U1/n995 ) );
  AO22_X0P5M_A12TL \U1/U981  ( .A0(\U1/n1104 ), .A1(\U1/key [37]), .B0(\U1/n1 ), .B1(Kin[37]), .Y(\U1/n994 ) );
  AO22_X0P5M_A12TL \U1/U980  ( .A0(\U1/n1107 ), .A1(\U1/key [36]), .B0(\U1/n1 ), .B1(Kin[36]), .Y(\U1/n993 ) );
  AO22_X0P5M_A12TL \U1/U979  ( .A0(\U1/n1105 ), .A1(\U1/key [35]), .B0(\U1/n1 ), .B1(Kin[35]), .Y(\U1/n992 ) );
  AO22_X0P5M_A12TL \U1/U978  ( .A0(\U1/n1104 ), .A1(\U1/key [34]), .B0(\U1/n1 ), .B1(Kin[34]), .Y(\U1/n991 ) );
  AO22_X0P5M_A12TL \U1/U977  ( .A0(\U1/n1105 ), .A1(\U1/key [33]), .B0(\U1/n1 ), .B1(Kin[33]), .Y(\U1/n990 ) );
  AO22_X0P5M_A12TL \U1/U976  ( .A0(\U1/n1104 ), .A1(\U1/key [32]), .B0(\U1/n1 ), .B1(Kin[32]), .Y(\U1/n989 ) );
  AO22_X0P5M_A12TL \U1/U975  ( .A0(\U1/n1107 ), .A1(\U1/key [31]), .B0(\U1/n1 ), .B1(Kin[31]), .Y(\U1/n988 ) );
  AO22_X0P5M_A12TL \U1/U974  ( .A0(\U1/n1106 ), .A1(\U1/key [30]), .B0(\U1/n1 ), .B1(Kin[30]), .Y(\U1/n987 ) );
  AO22_X0P5M_A12TL \U1/U973  ( .A0(\U1/n1105 ), .A1(\U1/key [29]), .B0(\U1/n1 ), .B1(Kin[29]), .Y(\U1/n986 ) );
  AO22_X0P5M_A12TL \U1/U972  ( .A0(\U1/n1104 ), .A1(\U1/key [28]), .B0(\U1/n1 ), .B1(Kin[28]), .Y(\U1/n985 ) );
  AO22_X0P5M_A12TL \U1/U971  ( .A0(\U1/n1107 ), .A1(\U1/key [27]), .B0(\U1/n1 ), .B1(Kin[27]), .Y(\U1/n984 ) );
  AO22_X0P5M_A12TL \U1/U970  ( .A0(\U1/n1106 ), .A1(\U1/key [26]), .B0(\U1/n1 ), .B1(Kin[26]), .Y(\U1/n983 ) );
  AO22_X0P5M_A12TL \U1/U969  ( .A0(\U1/n1105 ), .A1(\U1/key [25]), .B0(\U1/n1 ), .B1(Kin[25]), .Y(\U1/n982 ) );
  AO22_X0P5M_A12TL \U1/U968  ( .A0(\U1/n1104 ), .A1(\U1/key [24]), .B0(\U1/n1 ), .B1(Kin[24]), .Y(\U1/n981 ) );
  AO22_X0P5M_A12TL \U1/U967  ( .A0(\U1/n1105 ), .A1(\U1/key [23]), .B0(\U1/n1 ), .B1(Kin[23]), .Y(\U1/n980 ) );
  AO22_X0P5M_A12TL \U1/U966  ( .A0(\U1/n1105 ), .A1(\U1/key [22]), .B0(\U1/n1 ), .B1(Kin[22]), .Y(\U1/n979 ) );
  AO22_X0P5M_A12TL \U1/U965  ( .A0(\U1/n1105 ), .A1(\U1/key [21]), .B0(\U1/n1 ), .B1(Kin[21]), .Y(\U1/n978 ) );
  AO22_X0P5M_A12TL \U1/U964  ( .A0(\U1/n1105 ), .A1(\U1/key [20]), .B0(\U1/n1 ), .B1(Kin[20]), .Y(\U1/n977 ) );
  AO22_X0P5M_A12TL \U1/U963  ( .A0(\U1/n1105 ), .A1(\U1/key [19]), .B0(\U1/n1 ), .B1(Kin[19]), .Y(\U1/n976 ) );
  AO22_X0P5M_A12TL \U1/U962  ( .A0(\U1/n1105 ), .A1(\U1/key [18]), .B0(\U1/n1 ), .B1(Kin[18]), .Y(\U1/n975 ) );
  AO22_X0P5M_A12TL \U1/U961  ( .A0(\U1/n1105 ), .A1(\U1/key [17]), .B0(\U1/n1 ), .B1(Kin[17]), .Y(\U1/n974 ) );
  AO22_X0P5M_A12TL \U1/U960  ( .A0(\U1/n1105 ), .A1(\U1/key [16]), .B0(\U1/n1 ), .B1(Kin[16]), .Y(\U1/n973 ) );
  AO22_X0P5M_A12TL \U1/U959  ( .A0(\U1/n1105 ), .A1(\U1/key [15]), .B0(\U1/n1 ), .B1(Kin[15]), .Y(\U1/n972 ) );
  AO22_X0P5M_A12TL \U1/U958  ( .A0(\U1/n1105 ), .A1(\U1/key [14]), .B0(
        \U1/n1108 ), .B1(Kin[14]), .Y(\U1/n971 ) );
  AO22_X0P5M_A12TL \U1/U957  ( .A0(\U1/n1105 ), .A1(\U1/key [13]), .B0(
        \U1/n1108 ), .B1(Kin[13]), .Y(\U1/n970 ) );
  AO22_X0P5M_A12TL \U1/U956  ( .A0(\U1/n1105 ), .A1(\U1/key [12]), .B0(
        \U1/n1108 ), .B1(Kin[12]), .Y(\U1/n969 ) );
  AO22_X0P5M_A12TL \U1/U955  ( .A0(\U1/n1104 ), .A1(\U1/key [11]), .B0(
        \U1/n1108 ), .B1(Kin[11]), .Y(\U1/n968 ) );
  AO22_X0P5M_A12TL \U1/U954  ( .A0(\U1/n1104 ), .A1(\U1/key [10]), .B0(
        \U1/n1108 ), .B1(Kin[10]), .Y(\U1/n967 ) );
  AO22_X0P5M_A12TL \U1/U953  ( .A0(\U1/n1104 ), .A1(\U1/key [9]), .B0(
        \U1/n1108 ), .B1(Kin[9]), .Y(\U1/n966 ) );
  AO22_X0P5M_A12TL \U1/U952  ( .A0(\U1/n1104 ), .A1(\U1/key [8]), .B0(
        \U1/n1108 ), .B1(Kin[8]), .Y(\U1/n965 ) );
  AO22_X0P5M_A12TL \U1/U951  ( .A0(\U1/n1104 ), .A1(\U1/key [7]), .B0(
        \U1/n1108 ), .B1(Kin[7]), .Y(\U1/n964 ) );
  AO22_X0P5M_A12TL \U1/U950  ( .A0(\U1/n1104 ), .A1(\U1/key [6]), .B0(
        \U1/n1108 ), .B1(Kin[6]), .Y(\U1/n963 ) );
  AO22_X0P5M_A12TL \U1/U949  ( .A0(\U1/n1104 ), .A1(\U1/key [5]), .B0(
        \U1/n1108 ), .B1(Kin[5]), .Y(\U1/n962 ) );
  AO22_X0P5M_A12TL \U1/U948  ( .A0(\U1/n1104 ), .A1(\U1/key [4]), .B0(
        \U1/n1108 ), .B1(Kin[4]), .Y(\U1/n961 ) );
  AO22_X0P5M_A12TL \U1/U947  ( .A0(\U1/n1104 ), .A1(\U1/key [3]), .B0(
        \U1/n1108 ), .B1(Kin[3]), .Y(\U1/n960 ) );
  AO22_X0P5M_A12TL \U1/U946  ( .A0(\U1/n1104 ), .A1(\U1/key [2]), .B0(\U1/n1 ), 
        .B1(Kin[2]), .Y(\U1/n959 ) );
  AO22_X0P5M_A12TL \U1/U945  ( .A0(\U1/n1104 ), .A1(\U1/key [1]), .B0(\U1/n1 ), 
        .B1(Kin[1]), .Y(\U1/n958 ) );
  AO22_X0P5M_A12TL \U1/U944  ( .A0(\U1/n1104 ), .A1(\U1/key [0]), .B0(
        \U1/n1108 ), .B1(Kin[0]), .Y(\U1/n957 ) );
  NOR2_X0P5A_A12TL \U1/U943  ( .A(KDrdy2), .B(\U1/rnd [0]), .Y(\U1/n662 ) );
  AOI21B_X0P5M_A12TL \U1/U942  ( .A0(EN), .A1(\U1/n662 ), .B0N(\U1/n661 ), .Y(
        \U1/n669 ) );
  INV_X0P5B_A12TL \U1/U941  ( .A(\U1/n669 ), .Y(\U1/n663 ) );
  NAND2_X0P5A_A12TL \U1/U940  ( .A(\U1/n662 ), .B(\U1/n663 ), .Y(\U1/n665 ) );
  INV_X0P5B_A12TL \U1/U939  ( .A(\U1/rcon [7]), .Y(\U1/n664 ) );
  INV_X0P5B_A12TL \U1/U938  ( .A(KDrdy2), .Y(\U1/n659 ) );
  OAI222_X0P5M_A12TL \U1/U937  ( .A0(\U1/n808 ), .A1(\U1/n663 ), .B0(\U1/n665 ), .B1(\U1/n664 ), .C0(\U1/n669 ), .C1(\U1/n659 ), .Y(\U1/n956 ) );
  XNOR2_X0P5M_A12TL \U1/U936  ( .A(\U1/n664 ), .B(\U1/n808 ), .Y(\U1/n668 ) );
  OAI22_X0P5M_A12TL \U1/U935  ( .A0(\U1/n807 ), .A1(\U1/n663 ), .B0(\U1/n665 ), 
        .B1(\U1/n668 ), .Y(\U1/n955 ) );
  OAI22_X0P5M_A12TL \U1/U934  ( .A0(\U1/n806 ), .A1(\U1/n663 ), .B0(\U1/n807 ), 
        .B1(\U1/n665 ), .Y(\U1/n954 ) );
  XNOR2_X0P5M_A12TL \U1/U933  ( .A(\U1/n664 ), .B(\U1/n806 ), .Y(\U1/n667 ) );
  OAI22_X0P5M_A12TL \U1/U932  ( .A0(\U1/n805 ), .A1(\U1/n663 ), .B0(\U1/n665 ), 
        .B1(\U1/n667 ), .Y(\U1/n953 ) );
  XNOR2_X0P5M_A12TL \U1/U931  ( .A(\U1/n664 ), .B(\U1/n805 ), .Y(\U1/n666 ) );
  OAI22_X0P5M_A12TL \U1/U930  ( .A0(\U1/n804 ), .A1(\U1/n663 ), .B0(\U1/n665 ), 
        .B1(\U1/n666 ), .Y(\U1/n952 ) );
  OAI22_X0P5M_A12TL \U1/U929  ( .A0(\U1/n803 ), .A1(\U1/n663 ), .B0(\U1/n804 ), 
        .B1(\U1/n665 ), .Y(\U1/n951 ) );
  OAI22_X0P5M_A12TL \U1/U928  ( .A0(\U1/n802 ), .A1(\U1/n663 ), .B0(\U1/n803 ), 
        .B1(\U1/n665 ), .Y(\U1/n950 ) );
  OAI22_X0P5M_A12TL \U1/U927  ( .A0(\U1/n663 ), .A1(\U1/n664 ), .B0(\U1/n802 ), 
        .B1(\U1/n665 ), .Y(\U1/n949 ) );
  OAI21_X0P5M_A12TL \U1/U926  ( .A0(\U1/sel ), .A1(\U1/n662 ), .B0(EN), .Y(
        \U1/n660 ) );
  AND2_X0P5M_A12TL \U1/U925  ( .A(\U1/n660 ), .B(\U1/n661 ), .Y(\U1/n400 ) );
  NOR2_X0P5A_A12TL \U1/U924  ( .A(\U1/n659 ), .B(\U1/n400 ), .Y(\U1/n402 ) );
  XOR2_X0P5M_A12TL \U1/U923  ( .A(\U1/key [0]), .B(Din[0]), .Y(\U1/n658 ) );
  AOI22_X0P5M_A12TL \U1/U921  ( .A0(\U1/n1097 ), .A1(\U1/n658 ), .B0(
        \U1/dat_next [0]), .B1(\U1/n670 ), .Y(\U1/n657 ) );
  AO1B2_X0P5M_A12TL \U1/U920  ( .B0(Dout[0]), .B1(\U1/n1098 ), .A0N(\U1/n657 ), 
        .Y(\U1/n948 ) );
  XOR2_X0P5M_A12TL \U1/U919  ( .A(\U1/key [1]), .B(Din[1]), .Y(\U1/n656 ) );
  AOI22_X0P5M_A12TL \U1/U918  ( .A0(\U1/n1097 ), .A1(\U1/n656 ), .B0(
        \U1/dat_next [1]), .B1(\U1/n670 ), .Y(\U1/n655 ) );
  AO1B2_X0P5M_A12TL \U1/U917  ( .B0(Dout[1]), .B1(\U1/n1098 ), .A0N(\U1/n655 ), 
        .Y(\U1/n947 ) );
  XOR2_X0P5M_A12TL \U1/U916  ( .A(\U1/key [2]), .B(Din[2]), .Y(\U1/n654 ) );
  AOI22_X0P5M_A12TL \U1/U915  ( .A0(\U1/n1097 ), .A1(\U1/n654 ), .B0(
        \U1/dat_next [2]), .B1(\U1/n670 ), .Y(\U1/n653 ) );
  AO1B2_X0P5M_A12TL \U1/U914  ( .B0(Dout[2]), .B1(\U1/n1098 ), .A0N(\U1/n653 ), 
        .Y(\U1/n946 ) );
  XOR2_X0P5M_A12TL \U1/U913  ( .A(\U1/key [3]), .B(Din[3]), .Y(\U1/n652 ) );
  AOI22_X0P5M_A12TL \U1/U912  ( .A0(\U1/n1097 ), .A1(\U1/n652 ), .B0(
        \U1/dat_next [3]), .B1(\U1/n670 ), .Y(\U1/n651 ) );
  AO1B2_X0P5M_A12TL \U1/U911  ( .B0(Dout[3]), .B1(\U1/n1098 ), .A0N(\U1/n651 ), 
        .Y(\U1/n945 ) );
  XOR2_X0P5M_A12TL \U1/U910  ( .A(\U1/key [4]), .B(Din[4]), .Y(\U1/n650 ) );
  AOI22_X0P5M_A12TL \U1/U909  ( .A0(\U1/n1097 ), .A1(\U1/n650 ), .B0(
        \U1/dat_next [4]), .B1(\U1/n670 ), .Y(\U1/n649 ) );
  AO1B2_X0P5M_A12TL \U1/U908  ( .B0(Dout[4]), .B1(\U1/n1098 ), .A0N(\U1/n649 ), 
        .Y(\U1/n944 ) );
  XOR2_X0P5M_A12TL \U1/U907  ( .A(\U1/key [5]), .B(Din[5]), .Y(\U1/n648 ) );
  AOI22_X0P5M_A12TL \U1/U906  ( .A0(\U1/n1097 ), .A1(\U1/n648 ), .B0(
        \U1/dat_next [5]), .B1(\U1/n670 ), .Y(\U1/n647 ) );
  AO1B2_X0P5M_A12TL \U1/U905  ( .B0(Dout[5]), .B1(\U1/n1098 ), .A0N(\U1/n647 ), 
        .Y(\U1/n943 ) );
  XOR2_X0P5M_A12TL \U1/U904  ( .A(\U1/key [6]), .B(Din[6]), .Y(\U1/n646 ) );
  AOI22_X0P5M_A12TL \U1/U903  ( .A0(\U1/n1097 ), .A1(\U1/n646 ), .B0(
        \U1/dat_next [6]), .B1(\U1/n670 ), .Y(\U1/n645 ) );
  AO1B2_X0P5M_A12TL \U1/U902  ( .B0(Dout[6]), .B1(\U1/n1098 ), .A0N(\U1/n645 ), 
        .Y(\U1/n942 ) );
  XOR2_X0P5M_A12TL \U1/U901  ( .A(\U1/key [7]), .B(Din[7]), .Y(\U1/n644 ) );
  AOI22_X0P5M_A12TL \U1/U900  ( .A0(\U1/n1097 ), .A1(\U1/n644 ), .B0(
        \U1/dat_next [7]), .B1(\U1/n670 ), .Y(\U1/n643 ) );
  AO1B2_X0P5M_A12TL \U1/U899  ( .B0(Dout[7]), .B1(\U1/n1098 ), .A0N(\U1/n643 ), 
        .Y(\U1/n941 ) );
  XOR2_X0P5M_A12TL \U1/U898  ( .A(\U1/key [8]), .B(Din[8]), .Y(\U1/n642 ) );
  AOI22_X0P5M_A12TL \U1/U897  ( .A0(\U1/n1097 ), .A1(\U1/n642 ), .B0(
        \U1/dat_next [8]), .B1(\U1/n670 ), .Y(\U1/n641 ) );
  AO1B2_X0P5M_A12TL \U1/U896  ( .B0(Dout[8]), .B1(\U1/n1098 ), .A0N(\U1/n641 ), 
        .Y(\U1/n940 ) );
  XOR2_X0P5M_A12TL \U1/U895  ( .A(\U1/key [9]), .B(Din[9]), .Y(\U1/n640 ) );
  AOI22_X0P5M_A12TL \U1/U894  ( .A0(\U1/n1097 ), .A1(\U1/n640 ), .B0(
        \U1/dat_next [9]), .B1(\U1/n670 ), .Y(\U1/n639 ) );
  AO1B2_X0P5M_A12TL \U1/U893  ( .B0(Dout[9]), .B1(\U1/n1098 ), .A0N(\U1/n639 ), 
        .Y(\U1/n939 ) );
  XOR2_X0P5M_A12TL \U1/U892  ( .A(\U1/key [10]), .B(Din[10]), .Y(\U1/n638 ) );
  AOI22_X0P5M_A12TL \U1/U891  ( .A0(\U1/n1097 ), .A1(\U1/n638 ), .B0(
        \U1/dat_next [10]), .B1(\U1/n670 ), .Y(\U1/n637 ) );
  AO1B2_X0P5M_A12TL \U1/U890  ( .B0(Dout[10]), .B1(\U1/n1098 ), .A0N(\U1/n637 ), .Y(\U1/n938 ) );
  XOR2_X0P5M_A12TL \U1/U889  ( .A(\U1/key [11]), .B(Din[11]), .Y(\U1/n636 ) );
  AOI22_X0P5M_A12TL \U1/U888  ( .A0(\U1/n1097 ), .A1(\U1/n636 ), .B0(
        \U1/dat_next [11]), .B1(\U1/n670 ), .Y(\U1/n635 ) );
  AO1B2_X0P5M_A12TL \U1/U887  ( .B0(Dout[11]), .B1(\U1/n1098 ), .A0N(\U1/n635 ), .Y(\U1/n937 ) );
  XOR2_X0P5M_A12TL \U1/U886  ( .A(\U1/key [12]), .B(Din[12]), .Y(\U1/n634 ) );
  AOI22_X0P5M_A12TL \U1/U885  ( .A0(\U1/n1097 ), .A1(\U1/n634 ), .B0(
        \U1/dat_next [12]), .B1(\U1/n670 ), .Y(\U1/n633 ) );
  AO1B2_X0P5M_A12TL \U1/U884  ( .B0(Dout[12]), .B1(\U1/n1098 ), .A0N(\U1/n633 ), .Y(\U1/n936 ) );
  XOR2_X0P5M_A12TL \U1/U883  ( .A(\U1/key [13]), .B(Din[13]), .Y(\U1/n632 ) );
  AOI22_X0P5M_A12TL \U1/U882  ( .A0(\U1/n1096 ), .A1(\U1/n632 ), .B0(
        \U1/dat_next [13]), .B1(\U1/n670 ), .Y(\U1/n631 ) );
  AO1B2_X0P5M_A12TL \U1/U881  ( .B0(Dout[13]), .B1(\U1/n1098 ), .A0N(\U1/n631 ), .Y(\U1/n935 ) );
  XOR2_X0P5M_A12TL \U1/U880  ( .A(\U1/key [14]), .B(Din[14]), .Y(\U1/n630 ) );
  AOI22_X0P5M_A12TL \U1/U879  ( .A0(\U1/n1095 ), .A1(\U1/n630 ), .B0(
        \U1/dat_next [14]), .B1(\U1/n670 ), .Y(\U1/n629 ) );
  AO1B2_X0P5M_A12TL \U1/U878  ( .B0(Dout[14]), .B1(\U1/n1098 ), .A0N(\U1/n629 ), .Y(\U1/n934 ) );
  XOR2_X0P5M_A12TL \U1/U877  ( .A(\U1/key [15]), .B(Din[15]), .Y(\U1/n628 ) );
  AOI22_X0P5M_A12TL \U1/U876  ( .A0(\U1/n1097 ), .A1(\U1/n628 ), .B0(
        \U1/dat_next [15]), .B1(\U1/n670 ), .Y(\U1/n627 ) );
  AO1B2_X0P5M_A12TL \U1/U875  ( .B0(Dout[15]), .B1(\U1/n1098 ), .A0N(\U1/n627 ), .Y(\U1/n933 ) );
  XOR2_X0P5M_A12TL \U1/U874  ( .A(\U1/key [16]), .B(Din[16]), .Y(\U1/n626 ) );
  AOI22_X0P5M_A12TL \U1/U873  ( .A0(\U1/n1097 ), .A1(\U1/n626 ), .B0(
        \U1/dat_next [16]), .B1(\U1/n670 ), .Y(\U1/n625 ) );
  AO1B2_X0P5M_A12TL \U1/U872  ( .B0(Dout[16]), .B1(\U1/n1098 ), .A0N(\U1/n625 ), .Y(\U1/n932 ) );
  XOR2_X0P5M_A12TL \U1/U871  ( .A(\U1/key [17]), .B(Din[17]), .Y(\U1/n624 ) );
  AOI22_X0P5M_A12TL \U1/U870  ( .A0(\U1/n1097 ), .A1(\U1/n624 ), .B0(
        \U1/dat_next [17]), .B1(\U1/n670 ), .Y(\U1/n623 ) );
  AO1B2_X0P5M_A12TL \U1/U869  ( .B0(Dout[17]), .B1(\U1/n1098 ), .A0N(\U1/n623 ), .Y(\U1/n931 ) );
  XOR2_X0P5M_A12TL \U1/U868  ( .A(\U1/key [18]), .B(Din[18]), .Y(\U1/n622 ) );
  AOI22_X0P5M_A12TL \U1/U867  ( .A0(\U1/n1097 ), .A1(\U1/n622 ), .B0(
        \U1/dat_next [18]), .B1(\U1/n670 ), .Y(\U1/n621 ) );
  AO1B2_X0P5M_A12TL \U1/U866  ( .B0(Dout[18]), .B1(\U1/n1098 ), .A0N(\U1/n621 ), .Y(\U1/n930 ) );
  XOR2_X0P5M_A12TL \U1/U865  ( .A(\U1/key [19]), .B(Din[19]), .Y(\U1/n620 ) );
  AOI22_X0P5M_A12TL \U1/U864  ( .A0(\U1/n1097 ), .A1(\U1/n620 ), .B0(
        \U1/dat_next [19]), .B1(\U1/n670 ), .Y(\U1/n619 ) );
  AO1B2_X0P5M_A12TL \U1/U863  ( .B0(Dout[19]), .B1(\U1/n1098 ), .A0N(\U1/n619 ), .Y(\U1/n929 ) );
  XOR2_X0P5M_A12TL \U1/U862  ( .A(\U1/key [20]), .B(Din[20]), .Y(\U1/n618 ) );
  AOI22_X0P5M_A12TL \U1/U861  ( .A0(\U1/n1097 ), .A1(\U1/n618 ), .B0(
        \U1/dat_next [20]), .B1(\U1/n670 ), .Y(\U1/n617 ) );
  AO1B2_X0P5M_A12TL \U1/U860  ( .B0(Dout[20]), .B1(\U1/n1098 ), .A0N(\U1/n617 ), .Y(\U1/n928 ) );
  XOR2_X0P5M_A12TL \U1/U859  ( .A(\U1/key [21]), .B(Din[21]), .Y(\U1/n616 ) );
  AOI22_X0P5M_A12TL \U1/U858  ( .A0(\U1/n1097 ), .A1(\U1/n616 ), .B0(
        \U1/dat_next [21]), .B1(\U1/n670 ), .Y(\U1/n615 ) );
  AO1B2_X0P5M_A12TL \U1/U857  ( .B0(Dout[21]), .B1(\U1/n1098 ), .A0N(\U1/n615 ), .Y(\U1/n927 ) );
  XOR2_X0P5M_A12TL \U1/U856  ( .A(\U1/key [22]), .B(Din[22]), .Y(\U1/n614 ) );
  AOI22_X0P5M_A12TL \U1/U855  ( .A0(\U1/n1097 ), .A1(\U1/n614 ), .B0(
        \U1/dat_next [22]), .B1(\U1/n670 ), .Y(\U1/n613 ) );
  AO1B2_X0P5M_A12TL \U1/U854  ( .B0(Dout[22]), .B1(\U1/n1098 ), .A0N(\U1/n613 ), .Y(\U1/n926 ) );
  XOR2_X0P5M_A12TL \U1/U853  ( .A(\U1/key [23]), .B(Din[23]), .Y(\U1/n612 ) );
  AOI22_X0P5M_A12TL \U1/U852  ( .A0(\U1/n1097 ), .A1(\U1/n612 ), .B0(
        \U1/dat_next [23]), .B1(\U1/n670 ), .Y(\U1/n611 ) );
  AO1B2_X0P5M_A12TL \U1/U851  ( .B0(Dout[23]), .B1(\U1/n1098 ), .A0N(\U1/n611 ), .Y(\U1/n925 ) );
  XOR2_X0P5M_A12TL \U1/U850  ( .A(\U1/key [24]), .B(Din[24]), .Y(\U1/n610 ) );
  AOI22_X0P5M_A12TL \U1/U849  ( .A0(\U1/n1097 ), .A1(\U1/n610 ), .B0(
        \U1/dat_next [24]), .B1(\U1/n670 ), .Y(\U1/n609 ) );
  AO1B2_X0P5M_A12TL \U1/U848  ( .B0(Dout[24]), .B1(\U1/n1098 ), .A0N(\U1/n609 ), .Y(\U1/n924 ) );
  XOR2_X0P5M_A12TL \U1/U847  ( .A(\U1/key [25]), .B(Din[25]), .Y(\U1/n608 ) );
  AOI22_X0P5M_A12TL \U1/U846  ( .A0(\U1/n1097 ), .A1(\U1/n608 ), .B0(
        \U1/dat_next [25]), .B1(\U1/n670 ), .Y(\U1/n607 ) );
  AO1B2_X0P5M_A12TL \U1/U845  ( .B0(Dout[25]), .B1(\U1/n1098 ), .A0N(\U1/n607 ), .Y(\U1/n923 ) );
  XOR2_X0P5M_A12TL \U1/U844  ( .A(\U1/key [26]), .B(Din[26]), .Y(\U1/n606 ) );
  AOI22_X0P5M_A12TL \U1/U843  ( .A0(\U1/n1095 ), .A1(\U1/n606 ), .B0(
        \U1/dat_next [26]), .B1(\U1/n404 ), .Y(\U1/n605 ) );
  AO1B2_X0P5M_A12TL \U1/U842  ( .B0(Dout[26]), .B1(\U1/n1098 ), .A0N(\U1/n605 ), .Y(\U1/n922 ) );
  XOR2_X0P5M_A12TL \U1/U841  ( .A(\U1/key [27]), .B(Din[27]), .Y(\U1/n604 ) );
  AOI22_X0P5M_A12TL \U1/U840  ( .A0(\U1/n1095 ), .A1(\U1/n604 ), .B0(
        \U1/dat_next [27]), .B1(\U1/n404 ), .Y(\U1/n603 ) );
  AO1B2_X0P5M_A12TL \U1/U839  ( .B0(Dout[27]), .B1(\U1/n1098 ), .A0N(\U1/n603 ), .Y(\U1/n921 ) );
  XOR2_X0P5M_A12TL \U1/U838  ( .A(\U1/key [28]), .B(Din[28]), .Y(\U1/n602 ) );
  AOI22_X0P5M_A12TL \U1/U837  ( .A0(\U1/n1095 ), .A1(\U1/n602 ), .B0(
        \U1/dat_next [28]), .B1(\U1/n404 ), .Y(\U1/n601 ) );
  AO1B2_X0P5M_A12TL \U1/U836  ( .B0(Dout[28]), .B1(\U1/n1098 ), .A0N(\U1/n601 ), .Y(\U1/n920 ) );
  XOR2_X0P5M_A12TL \U1/U835  ( .A(\U1/key [29]), .B(Din[29]), .Y(\U1/n600 ) );
  AOI22_X0P5M_A12TL \U1/U834  ( .A0(\U1/n1095 ), .A1(\U1/n600 ), .B0(
        \U1/dat_next [29]), .B1(\U1/n404 ), .Y(\U1/n599 ) );
  AO1B2_X0P5M_A12TL \U1/U833  ( .B0(Dout[29]), .B1(\U1/n1098 ), .A0N(\U1/n599 ), .Y(\U1/n919 ) );
  XOR2_X0P5M_A12TL \U1/U832  ( .A(\U1/key [30]), .B(Din[30]), .Y(\U1/n598 ) );
  AOI22_X0P5M_A12TL \U1/U831  ( .A0(\U1/n1095 ), .A1(\U1/n598 ), .B0(
        \U1/dat_next [30]), .B1(\U1/n670 ), .Y(\U1/n597 ) );
  AO1B2_X0P5M_A12TL \U1/U830  ( .B0(Dout[30]), .B1(\U1/n1098 ), .A0N(\U1/n597 ), .Y(\U1/n918 ) );
  XOR2_X0P5M_A12TL \U1/U829  ( .A(\U1/key [31]), .B(Din[31]), .Y(\U1/n596 ) );
  AOI22_X0P5M_A12TL \U1/U828  ( .A0(\U1/n1095 ), .A1(\U1/n596 ), .B0(
        \U1/dat_next [31]), .B1(\U1/n670 ), .Y(\U1/n595 ) );
  AO1B2_X0P5M_A12TL \U1/U827  ( .B0(Dout[31]), .B1(\U1/n1098 ), .A0N(\U1/n595 ), .Y(\U1/n917 ) );
  XOR2_X0P5M_A12TL \U1/U826  ( .A(\U1/key [32]), .B(Din[32]), .Y(\U1/n594 ) );
  AOI22_X0P5M_A12TL \U1/U825  ( .A0(\U1/n1095 ), .A1(\U1/n594 ), .B0(
        \U1/dat_next [32]), .B1(\U1/n670 ), .Y(\U1/n593 ) );
  AO1B2_X0P5M_A12TL \U1/U824  ( .B0(Dout[32]), .B1(\U1/n1098 ), .A0N(\U1/n593 ), .Y(\U1/n916 ) );
  XOR2_X0P5M_A12TL \U1/U823  ( .A(\U1/key [33]), .B(Din[33]), .Y(\U1/n592 ) );
  AOI22_X0P5M_A12TL \U1/U822  ( .A0(\U1/n1095 ), .A1(\U1/n592 ), .B0(
        \U1/dat_next [33]), .B1(\U1/n670 ), .Y(\U1/n591 ) );
  AO1B2_X0P5M_A12TL \U1/U821  ( .B0(Dout[33]), .B1(\U1/n1098 ), .A0N(\U1/n591 ), .Y(\U1/n915 ) );
  XOR2_X0P5M_A12TL \U1/U820  ( .A(\U1/key [34]), .B(Din[34]), .Y(\U1/n590 ) );
  AOI22_X0P5M_A12TL \U1/U819  ( .A0(\U1/n1095 ), .A1(\U1/n590 ), .B0(
        \U1/dat_next [34]), .B1(\U1/n670 ), .Y(\U1/n589 ) );
  AO1B2_X0P5M_A12TL \U1/U818  ( .B0(Dout[34]), .B1(\U1/n1098 ), .A0N(\U1/n589 ), .Y(\U1/n914 ) );
  XOR2_X0P5M_A12TL \U1/U817  ( .A(\U1/key [35]), .B(Din[35]), .Y(\U1/n588 ) );
  AOI22_X0P5M_A12TL \U1/U816  ( .A0(\U1/n1095 ), .A1(\U1/n588 ), .B0(
        \U1/dat_next [35]), .B1(\U1/n670 ), .Y(\U1/n587 ) );
  AO1B2_X0P5M_A12TL \U1/U815  ( .B0(Dout[35]), .B1(\U1/n1098 ), .A0N(\U1/n587 ), .Y(\U1/n913 ) );
  XOR2_X0P5M_A12TL \U1/U814  ( .A(\U1/key [36]), .B(Din[36]), .Y(\U1/n586 ) );
  AOI22_X0P5M_A12TL \U1/U813  ( .A0(\U1/n1095 ), .A1(\U1/n586 ), .B0(
        \U1/dat_next [36]), .B1(\U1/n670 ), .Y(\U1/n585 ) );
  AO1B2_X0P5M_A12TL \U1/U812  ( .B0(Dout[36]), .B1(\U1/n1098 ), .A0N(\U1/n585 ), .Y(\U1/n912 ) );
  XOR2_X0P5M_A12TL \U1/U811  ( .A(\U1/key [37]), .B(Din[37]), .Y(\U1/n584 ) );
  AOI22_X0P5M_A12TL \U1/U810  ( .A0(\U1/n1095 ), .A1(\U1/n584 ), .B0(
        \U1/dat_next [37]), .B1(\U1/n670 ), .Y(\U1/n583 ) );
  AO1B2_X0P5M_A12TL \U1/U809  ( .B0(Dout[37]), .B1(\U1/n1098 ), .A0N(\U1/n583 ), .Y(\U1/n911 ) );
  XOR2_X0P5M_A12TL \U1/U808  ( .A(\U1/key [38]), .B(Din[38]), .Y(\U1/n582 ) );
  AOI22_X0P5M_A12TL \U1/U807  ( .A0(\U1/n1095 ), .A1(\U1/n582 ), .B0(
        \U1/dat_next [38]), .B1(\U1/n670 ), .Y(\U1/n581 ) );
  AO1B2_X0P5M_A12TL \U1/U806  ( .B0(Dout[38]), .B1(\U1/n1098 ), .A0N(\U1/n581 ), .Y(\U1/n910 ) );
  XOR2_X0P5M_A12TL \U1/U805  ( .A(\U1/key [39]), .B(Din[39]), .Y(\U1/n580 ) );
  AOI22_X0P5M_A12TL \U1/U804  ( .A0(\U1/n1096 ), .A1(\U1/n580 ), .B0(
        \U1/dat_next [39]), .B1(\U1/n670 ), .Y(\U1/n579 ) );
  AO1B2_X0P5M_A12TL \U1/U803  ( .B0(Dout[39]), .B1(\U1/n1098 ), .A0N(\U1/n579 ), .Y(\U1/n909 ) );
  XOR2_X0P5M_A12TL \U1/U802  ( .A(\U1/key [40]), .B(Din[40]), .Y(\U1/n578 ) );
  AOI22_X0P5M_A12TL \U1/U801  ( .A0(\U1/n1096 ), .A1(\U1/n578 ), .B0(
        \U1/dat_next [40]), .B1(\U1/n670 ), .Y(\U1/n577 ) );
  AO1B2_X0P5M_A12TL \U1/U800  ( .B0(Dout[40]), .B1(\U1/n1098 ), .A0N(\U1/n577 ), .Y(\U1/n908 ) );
  XOR2_X0P5M_A12TL \U1/U799  ( .A(\U1/key [41]), .B(Din[41]), .Y(\U1/n576 ) );
  AOI22_X0P5M_A12TL \U1/U798  ( .A0(\U1/n1096 ), .A1(\U1/n576 ), .B0(
        \U1/dat_next [41]), .B1(\U1/n670 ), .Y(\U1/n575 ) );
  AO1B2_X0P5M_A12TL \U1/U797  ( .B0(Dout[41]), .B1(\U1/n1098 ), .A0N(\U1/n575 ), .Y(\U1/n907 ) );
  XOR2_X0P5M_A12TL \U1/U796  ( .A(\U1/key [42]), .B(Din[42]), .Y(\U1/n574 ) );
  AOI22_X0P5M_A12TL \U1/U795  ( .A0(\U1/n1096 ), .A1(\U1/n574 ), .B0(
        \U1/dat_next [42]), .B1(\U1/n670 ), .Y(\U1/n573 ) );
  AO1B2_X0P5M_A12TL \U1/U794  ( .B0(Dout[42]), .B1(\U1/n1098 ), .A0N(\U1/n573 ), .Y(\U1/n906 ) );
  XOR2_X0P5M_A12TL \U1/U793  ( .A(\U1/key [43]), .B(Din[43]), .Y(\U1/n572 ) );
  AOI22_X0P5M_A12TL \U1/U792  ( .A0(\U1/n1096 ), .A1(\U1/n572 ), .B0(
        \U1/dat_next [43]), .B1(\U1/n670 ), .Y(\U1/n571 ) );
  AO1B2_X0P5M_A12TL \U1/U791  ( .B0(Dout[43]), .B1(\U1/n1098 ), .A0N(\U1/n571 ), .Y(\U1/n905 ) );
  XOR2_X0P5M_A12TL \U1/U790  ( .A(\U1/key [44]), .B(Din[44]), .Y(\U1/n570 ) );
  AOI22_X0P5M_A12TL \U1/U789  ( .A0(\U1/n1096 ), .A1(\U1/n570 ), .B0(
        \U1/dat_next [44]), .B1(\U1/n670 ), .Y(\U1/n569 ) );
  AO1B2_X0P5M_A12TL \U1/U788  ( .B0(Dout[44]), .B1(\U1/n1098 ), .A0N(\U1/n569 ), .Y(\U1/n904 ) );
  XOR2_X0P5M_A12TL \U1/U787  ( .A(\U1/key [45]), .B(Din[45]), .Y(\U1/n568 ) );
  AOI22_X0P5M_A12TL \U1/U786  ( .A0(\U1/n1096 ), .A1(\U1/n568 ), .B0(
        \U1/dat_next [45]), .B1(\U1/n670 ), .Y(\U1/n567 ) );
  AO1B2_X0P5M_A12TL \U1/U785  ( .B0(Dout[45]), .B1(\U1/n1098 ), .A0N(\U1/n567 ), .Y(\U1/n903 ) );
  XOR2_X0P5M_A12TL \U1/U784  ( .A(\U1/key [46]), .B(Din[46]), .Y(\U1/n566 ) );
  AOI22_X0P5M_A12TL \U1/U783  ( .A0(\U1/n1096 ), .A1(\U1/n566 ), .B0(
        \U1/dat_next [46]), .B1(\U1/n670 ), .Y(\U1/n565 ) );
  AO1B2_X0P5M_A12TL \U1/U782  ( .B0(Dout[46]), .B1(\U1/n1098 ), .A0N(\U1/n565 ), .Y(\U1/n902 ) );
  XOR2_X0P5M_A12TL \U1/U781  ( .A(\U1/key [47]), .B(Din[47]), .Y(\U1/n564 ) );
  AOI22_X0P5M_A12TL \U1/U780  ( .A0(\U1/n1096 ), .A1(\U1/n564 ), .B0(
        \U1/dat_next [47]), .B1(\U1/n670 ), .Y(\U1/n563 ) );
  AO1B2_X0P5M_A12TL \U1/U779  ( .B0(Dout[47]), .B1(\U1/n1098 ), .A0N(\U1/n563 ), .Y(\U1/n901 ) );
  XOR2_X0P5M_A12TL \U1/U778  ( .A(\U1/key [48]), .B(Din[48]), .Y(\U1/n562 ) );
  AOI22_X0P5M_A12TL \U1/U777  ( .A0(\U1/n1096 ), .A1(\U1/n562 ), .B0(
        \U1/dat_next [48]), .B1(\U1/n670 ), .Y(\U1/n561 ) );
  AO1B2_X0P5M_A12TL \U1/U776  ( .B0(Dout[48]), .B1(\U1/n1098 ), .A0N(\U1/n561 ), .Y(\U1/n900 ) );
  XOR2_X0P5M_A12TL \U1/U775  ( .A(\U1/key [49]), .B(Din[49]), .Y(\U1/n560 ) );
  AOI22_X0P5M_A12TL \U1/U774  ( .A0(\U1/n1096 ), .A1(\U1/n560 ), .B0(
        \U1/dat_next [49]), .B1(\U1/n670 ), .Y(\U1/n559 ) );
  AO1B2_X0P5M_A12TL \U1/U773  ( .B0(Dout[49]), .B1(\U1/n1098 ), .A0N(\U1/n559 ), .Y(\U1/n899 ) );
  XOR2_X0P5M_A12TL \U1/U772  ( .A(\U1/key [50]), .B(Din[50]), .Y(\U1/n558 ) );
  AOI22_X0P5M_A12TL \U1/U771  ( .A0(\U1/n1096 ), .A1(\U1/n558 ), .B0(
        \U1/dat_next [50]), .B1(\U1/n670 ), .Y(\U1/n557 ) );
  AO1B2_X0P5M_A12TL \U1/U770  ( .B0(Dout[50]), .B1(\U1/n1098 ), .A0N(\U1/n557 ), .Y(\U1/n898 ) );
  XOR2_X0P5M_A12TL \U1/U769  ( .A(\U1/key [51]), .B(Din[51]), .Y(\U1/n556 ) );
  AOI22_X0P5M_A12TL \U1/U768  ( .A0(\U1/n1096 ), .A1(\U1/n556 ), .B0(
        \U1/dat_next [51]), .B1(\U1/n670 ), .Y(\U1/n555 ) );
  AO1B2_X0P5M_A12TL \U1/U767  ( .B0(Dout[51]), .B1(\U1/n1098 ), .A0N(\U1/n555 ), .Y(\U1/n897 ) );
  XOR2_X0P5M_A12TL \U1/U766  ( .A(\U1/key [52]), .B(Din[52]), .Y(\U1/n554 ) );
  AOI22_X0P5M_A12TL \U1/U765  ( .A0(\U1/n402 ), .A1(\U1/n554 ), .B0(
        \U1/dat_next [52]), .B1(\U1/n670 ), .Y(\U1/n553 ) );
  AO1B2_X0P5M_A12TL \U1/U764  ( .B0(Dout[52]), .B1(\U1/n1098 ), .A0N(\U1/n553 ), .Y(\U1/n896 ) );
  XOR2_X0P5M_A12TL \U1/U763  ( .A(\U1/key [53]), .B(Din[53]), .Y(\U1/n552 ) );
  AOI22_X0P5M_A12TL \U1/U762  ( .A0(\U1/n1097 ), .A1(\U1/n552 ), .B0(
        \U1/dat_next [53]), .B1(\U1/n670 ), .Y(\U1/n551 ) );
  AO1B2_X0P5M_A12TL \U1/U761  ( .B0(Dout[53]), .B1(\U1/n1098 ), .A0N(\U1/n551 ), .Y(\U1/n895 ) );
  XOR2_X0P5M_A12TL \U1/U760  ( .A(\U1/key [54]), .B(Din[54]), .Y(\U1/n550 ) );
  AOI22_X0P5M_A12TL \U1/U759  ( .A0(\U1/n402 ), .A1(\U1/n550 ), .B0(
        \U1/dat_next [54]), .B1(\U1/n670 ), .Y(\U1/n549 ) );
  AO1B2_X0P5M_A12TL \U1/U758  ( .B0(Dout[54]), .B1(\U1/n1098 ), .A0N(\U1/n549 ), .Y(\U1/n894 ) );
  XOR2_X0P5M_A12TL \U1/U757  ( .A(\U1/key [55]), .B(Din[55]), .Y(\U1/n548 ) );
  AOI22_X0P5M_A12TL \U1/U756  ( .A0(\U1/n1097 ), .A1(\U1/n548 ), .B0(
        \U1/dat_next [55]), .B1(\U1/n670 ), .Y(\U1/n547 ) );
  AO1B2_X0P5M_A12TL \U1/U755  ( .B0(Dout[55]), .B1(\U1/n1098 ), .A0N(\U1/n547 ), .Y(\U1/n893 ) );
  XOR2_X0P5M_A12TL \U1/U754  ( .A(\U1/key [56]), .B(Din[56]), .Y(\U1/n546 ) );
  AOI22_X0P5M_A12TL \U1/U753  ( .A0(\U1/n402 ), .A1(\U1/n546 ), .B0(
        \U1/dat_next [56]), .B1(\U1/n670 ), .Y(\U1/n545 ) );
  AO1B2_X0P5M_A12TL \U1/U752  ( .B0(Dout[56]), .B1(\U1/n1098 ), .A0N(\U1/n545 ), .Y(\U1/n892 ) );
  XOR2_X0P5M_A12TL \U1/U751  ( .A(\U1/key [57]), .B(Din[57]), .Y(\U1/n544 ) );
  AOI22_X0P5M_A12TL \U1/U750  ( .A0(\U1/n1097 ), .A1(\U1/n544 ), .B0(
        \U1/dat_next [57]), .B1(\U1/n670 ), .Y(\U1/n543 ) );
  AO1B2_X0P5M_A12TL \U1/U749  ( .B0(Dout[57]), .B1(\U1/n1098 ), .A0N(\U1/n543 ), .Y(\U1/n891 ) );
  XOR2_X0P5M_A12TL \U1/U748  ( .A(\U1/key [58]), .B(Din[58]), .Y(\U1/n542 ) );
  AOI22_X0P5M_A12TL \U1/U747  ( .A0(\U1/n402 ), .A1(\U1/n542 ), .B0(
        \U1/dat_next [58]), .B1(\U1/n670 ), .Y(\U1/n541 ) );
  AO1B2_X0P5M_A12TL \U1/U746  ( .B0(Dout[58]), .B1(\U1/n1098 ), .A0N(\U1/n541 ), .Y(\U1/n890 ) );
  XOR2_X0P5M_A12TL \U1/U745  ( .A(\U1/key [59]), .B(Din[59]), .Y(\U1/n540 ) );
  AOI22_X0P5M_A12TL \U1/U744  ( .A0(\U1/n1097 ), .A1(\U1/n540 ), .B0(
        \U1/dat_next [59]), .B1(\U1/n670 ), .Y(\U1/n539 ) );
  AO1B2_X0P5M_A12TL \U1/U743  ( .B0(Dout[59]), .B1(\U1/n1098 ), .A0N(\U1/n539 ), .Y(\U1/n889 ) );
  XOR2_X0P5M_A12TL \U1/U742  ( .A(\U1/key [60]), .B(Din[60]), .Y(\U1/n538 ) );
  AOI22_X0P5M_A12TL \U1/U741  ( .A0(\U1/n402 ), .A1(\U1/n538 ), .B0(
        \U1/dat_next [60]), .B1(\U1/n670 ), .Y(\U1/n537 ) );
  AO1B2_X0P5M_A12TL \U1/U740  ( .B0(Dout[60]), .B1(\U1/n1098 ), .A0N(\U1/n537 ), .Y(\U1/n888 ) );
  XOR2_X0P5M_A12TL \U1/U739  ( .A(\U1/key [61]), .B(Din[61]), .Y(\U1/n536 ) );
  AOI22_X0P5M_A12TL \U1/U738  ( .A0(\U1/n1097 ), .A1(\U1/n536 ), .B0(
        \U1/dat_next [61]), .B1(\U1/n670 ), .Y(\U1/n535 ) );
  AO1B2_X0P5M_A12TL \U1/U737  ( .B0(Dout[61]), .B1(\U1/n1098 ), .A0N(\U1/n535 ), .Y(\U1/n887 ) );
  XOR2_X0P5M_A12TL \U1/U736  ( .A(\U1/key [62]), .B(Din[62]), .Y(\U1/n534 ) );
  AOI22_X0P5M_A12TL \U1/U735  ( .A0(\U1/n402 ), .A1(\U1/n534 ), .B0(
        \U1/dat_next [62]), .B1(\U1/n670 ), .Y(\U1/n533 ) );
  AO1B2_X0P5M_A12TL \U1/U734  ( .B0(Dout[62]), .B1(\U1/n1098 ), .A0N(\U1/n533 ), .Y(\U1/n886 ) );
  XOR2_X0P5M_A12TL \U1/U733  ( .A(\U1/key [63]), .B(Din[63]), .Y(\U1/n532 ) );
  AOI22_X0P5M_A12TL \U1/U732  ( .A0(\U1/n1097 ), .A1(\U1/n532 ), .B0(
        \U1/dat_next [63]), .B1(\U1/n670 ), .Y(\U1/n531 ) );
  AO1B2_X0P5M_A12TL \U1/U731  ( .B0(Dout[63]), .B1(\U1/n1098 ), .A0N(\U1/n531 ), .Y(\U1/n885 ) );
  XOR2_X0P5M_A12TL \U1/U730  ( .A(\U1/key [64]), .B(Din[64]), .Y(\U1/n530 ) );
  AOI22_X0P5M_A12TL \U1/U729  ( .A0(\U1/n1097 ), .A1(\U1/n530 ), .B0(
        \U1/dat_next [64]), .B1(\U1/n670 ), .Y(\U1/n529 ) );
  AO1B2_X0P5M_A12TL \U1/U728  ( .B0(Dout[64]), .B1(\U1/n1098 ), .A0N(\U1/n529 ), .Y(\U1/n884 ) );
  XOR2_X0P5M_A12TL \U1/U727  ( .A(\U1/key [65]), .B(Din[65]), .Y(\U1/n528 ) );
  AOI22_X0P5M_A12TL \U1/U726  ( .A0(\U1/n402 ), .A1(\U1/n528 ), .B0(
        \U1/dat_next [65]), .B1(\U1/n404 ), .Y(\U1/n527 ) );
  AO1B2_X0P5M_A12TL \U1/U725  ( .B0(Dout[65]), .B1(\U1/n1098 ), .A0N(\U1/n527 ), .Y(\U1/n883 ) );
  XOR2_X0P5M_A12TL \U1/U724  ( .A(\U1/key [66]), .B(Din[66]), .Y(\U1/n526 ) );
  AOI22_X0P5M_A12TL \U1/U723  ( .A0(\U1/n1097 ), .A1(\U1/n526 ), .B0(
        \U1/dat_next [66]), .B1(\U1/n404 ), .Y(\U1/n525 ) );
  AO1B2_X0P5M_A12TL \U1/U722  ( .B0(Dout[66]), .B1(\U1/n400 ), .A0N(\U1/n525 ), 
        .Y(\U1/n882 ) );
  XOR2_X0P5M_A12TL \U1/U721  ( .A(\U1/key [67]), .B(Din[67]), .Y(\U1/n524 ) );
  AOI22_X0P5M_A12TL \U1/U720  ( .A0(\U1/n1097 ), .A1(\U1/n524 ), .B0(
        \U1/dat_next [67]), .B1(\U1/n404 ), .Y(\U1/n523 ) );
  AO1B2_X0P5M_A12TL \U1/U719  ( .B0(Dout[67]), .B1(\U1/n400 ), .A0N(\U1/n523 ), 
        .Y(\U1/n881 ) );
  XOR2_X0P5M_A12TL \U1/U718  ( .A(\U1/key [68]), .B(Din[68]), .Y(\U1/n522 ) );
  AOI22_X0P5M_A12TL \U1/U717  ( .A0(\U1/n402 ), .A1(\U1/n522 ), .B0(
        \U1/dat_next [68]), .B1(\U1/n404 ), .Y(\U1/n521 ) );
  AO1B2_X0P5M_A12TL \U1/U716  ( .B0(Dout[68]), .B1(\U1/n400 ), .A0N(\U1/n521 ), 
        .Y(\U1/n880 ) );
  XOR2_X0P5M_A12TL \U1/U715  ( .A(\U1/key [69]), .B(Din[69]), .Y(\U1/n520 ) );
  AOI22_X0P5M_A12TL \U1/U714  ( .A0(\U1/n1097 ), .A1(\U1/n520 ), .B0(
        \U1/dat_next [69]), .B1(\U1/n404 ), .Y(\U1/n519 ) );
  AO1B2_X0P5M_A12TL \U1/U713  ( .B0(Dout[69]), .B1(\U1/n400 ), .A0N(\U1/n519 ), 
        .Y(\U1/n879 ) );
  XOR2_X0P5M_A12TL \U1/U712  ( .A(\U1/key [70]), .B(Din[70]), .Y(\U1/n518 ) );
  AOI22_X0P5M_A12TL \U1/U711  ( .A0(\U1/n1097 ), .A1(\U1/n518 ), .B0(
        \U1/dat_next [70]), .B1(\U1/n404 ), .Y(\U1/n517 ) );
  AO1B2_X0P5M_A12TL \U1/U710  ( .B0(Dout[70]), .B1(\U1/n400 ), .A0N(\U1/n517 ), 
        .Y(\U1/n878 ) );
  XOR2_X0P5M_A12TL \U1/U709  ( .A(\U1/key [71]), .B(Din[71]), .Y(\U1/n516 ) );
  AOI22_X0P5M_A12TL \U1/U708  ( .A0(\U1/n402 ), .A1(\U1/n516 ), .B0(
        \U1/dat_next [71]), .B1(\U1/n670 ), .Y(\U1/n515 ) );
  AO1B2_X0P5M_A12TL \U1/U707  ( .B0(Dout[71]), .B1(\U1/n400 ), .A0N(\U1/n515 ), 
        .Y(\U1/n877 ) );
  XOR2_X0P5M_A12TL \U1/U706  ( .A(\U1/key [72]), .B(Din[72]), .Y(\U1/n514 ) );
  AOI22_X0P5M_A12TL \U1/U705  ( .A0(\U1/n1097 ), .A1(\U1/n514 ), .B0(
        \U1/dat_next [72]), .B1(\U1/n404 ), .Y(\U1/n513 ) );
  AO1B2_X0P5M_A12TL \U1/U704  ( .B0(Dout[72]), .B1(\U1/n400 ), .A0N(\U1/n513 ), 
        .Y(\U1/n876 ) );
  XOR2_X0P5M_A12TL \U1/U703  ( .A(\U1/key [73]), .B(Din[73]), .Y(\U1/n512 ) );
  AOI22_X0P5M_A12TL \U1/U702  ( .A0(\U1/n402 ), .A1(\U1/n512 ), .B0(
        \U1/dat_next [73]), .B1(\U1/n670 ), .Y(\U1/n511 ) );
  AO1B2_X0P5M_A12TL \U1/U701  ( .B0(Dout[73]), .B1(\U1/n400 ), .A0N(\U1/n511 ), 
        .Y(\U1/n875 ) );
  XOR2_X0P5M_A12TL \U1/U700  ( .A(\U1/key [74]), .B(Din[74]), .Y(\U1/n510 ) );
  AOI22_X0P5M_A12TL \U1/U699  ( .A0(\U1/n1097 ), .A1(\U1/n510 ), .B0(
        \U1/dat_next [74]), .B1(\U1/n404 ), .Y(\U1/n509 ) );
  AO1B2_X0P5M_A12TL \U1/U698  ( .B0(Dout[74]), .B1(\U1/n400 ), .A0N(\U1/n509 ), 
        .Y(\U1/n874 ) );
  XOR2_X0P5M_A12TL \U1/U697  ( .A(\U1/key [75]), .B(Din[75]), .Y(\U1/n508 ) );
  AOI22_X0P5M_A12TL \U1/U696  ( .A0(\U1/n402 ), .A1(\U1/n508 ), .B0(
        \U1/dat_next [75]), .B1(\U1/n670 ), .Y(\U1/n507 ) );
  AO1B2_X0P5M_A12TL \U1/U695  ( .B0(Dout[75]), .B1(\U1/n400 ), .A0N(\U1/n507 ), 
        .Y(\U1/n873 ) );
  XOR2_X0P5M_A12TL \U1/U694  ( .A(\U1/key [76]), .B(Din[76]), .Y(\U1/n506 ) );
  AOI22_X0P5M_A12TL \U1/U693  ( .A0(\U1/n1097 ), .A1(\U1/n506 ), .B0(
        \U1/dat_next [76]), .B1(\U1/n404 ), .Y(\U1/n505 ) );
  AO1B2_X0P5M_A12TL \U1/U692  ( .B0(Dout[76]), .B1(\U1/n400 ), .A0N(\U1/n505 ), 
        .Y(\U1/n872 ) );
  XOR2_X0P5M_A12TL \U1/U691  ( .A(\U1/key [77]), .B(Din[77]), .Y(\U1/n504 ) );
  AOI22_X0P5M_A12TL \U1/U690  ( .A0(\U1/n1097 ), .A1(\U1/n504 ), .B0(
        \U1/dat_next [77]), .B1(\U1/n404 ), .Y(\U1/n503 ) );
  AO1B2_X0P5M_A12TL \U1/U689  ( .B0(Dout[77]), .B1(\U1/n400 ), .A0N(\U1/n503 ), 
        .Y(\U1/n871 ) );
  XOR2_X0P5M_A12TL \U1/U688  ( .A(\U1/key [78]), .B(Din[78]), .Y(\U1/n502 ) );
  AOI22_X0P5M_A12TL \U1/U687  ( .A0(\U1/n1097 ), .A1(\U1/n502 ), .B0(
        \U1/dat_next [78]), .B1(\U1/n404 ), .Y(\U1/n501 ) );
  AO1B2_X0P5M_A12TL \U1/U686  ( .B0(Dout[78]), .B1(\U1/n400 ), .A0N(\U1/n501 ), 
        .Y(\U1/n870 ) );
  XOR2_X0P5M_A12TL \U1/U685  ( .A(\U1/key [79]), .B(Din[79]), .Y(\U1/n500 ) );
  AOI22_X0P5M_A12TL \U1/U684  ( .A0(\U1/n1097 ), .A1(\U1/n500 ), .B0(
        \U1/dat_next [79]), .B1(\U1/n404 ), .Y(\U1/n499 ) );
  AO1B2_X0P5M_A12TL \U1/U683  ( .B0(Dout[79]), .B1(\U1/n400 ), .A0N(\U1/n499 ), 
        .Y(\U1/n869 ) );
  XOR2_X0P5M_A12TL \U1/U682  ( .A(\U1/key [80]), .B(Din[80]), .Y(\U1/n498 ) );
  AOI22_X0P5M_A12TL \U1/U681  ( .A0(\U1/n402 ), .A1(\U1/n498 ), .B0(
        \U1/dat_next [80]), .B1(\U1/n670 ), .Y(\U1/n497 ) );
  AO1B2_X0P5M_A12TL \U1/U680  ( .B0(Dout[80]), .B1(\U1/n400 ), .A0N(\U1/n497 ), 
        .Y(\U1/n868 ) );
  XOR2_X0P5M_A12TL \U1/U679  ( .A(\U1/key [81]), .B(Din[81]), .Y(\U1/n496 ) );
  AOI22_X0P5M_A12TL \U1/U678  ( .A0(\U1/n402 ), .A1(\U1/n496 ), .B0(
        \U1/dat_next [81]), .B1(\U1/n670 ), .Y(\U1/n495 ) );
  AO1B2_X0P5M_A12TL \U1/U677  ( .B0(Dout[81]), .B1(\U1/n400 ), .A0N(\U1/n495 ), 
        .Y(\U1/n867 ) );
  XOR2_X0P5M_A12TL \U1/U676  ( .A(\U1/key [82]), .B(Din[82]), .Y(\U1/n494 ) );
  AOI22_X0P5M_A12TL \U1/U675  ( .A0(\U1/n1097 ), .A1(\U1/n494 ), .B0(
        \U1/dat_next [82]), .B1(\U1/n670 ), .Y(\U1/n493 ) );
  AO1B2_X0P5M_A12TL \U1/U674  ( .B0(Dout[82]), .B1(\U1/n400 ), .A0N(\U1/n493 ), 
        .Y(\U1/n866 ) );
  XOR2_X0P5M_A12TL \U1/U673  ( .A(\U1/key [83]), .B(Din[83]), .Y(\U1/n492 ) );
  AOI22_X0P5M_A12TL \U1/U672  ( .A0(\U1/n1097 ), .A1(\U1/n492 ), .B0(
        \U1/dat_next [83]), .B1(\U1/n670 ), .Y(\U1/n491 ) );
  AO1B2_X0P5M_A12TL \U1/U671  ( .B0(Dout[83]), .B1(\U1/n400 ), .A0N(\U1/n491 ), 
        .Y(\U1/n865 ) );
  XOR2_X0P5M_A12TL \U1/U670  ( .A(\U1/key [84]), .B(Din[84]), .Y(\U1/n490 ) );
  AOI22_X0P5M_A12TL \U1/U669  ( .A0(\U1/n1097 ), .A1(\U1/n490 ), .B0(
        \U1/dat_next [84]), .B1(\U1/n404 ), .Y(\U1/n489 ) );
  AO1B2_X0P5M_A12TL \U1/U668  ( .B0(Dout[84]), .B1(\U1/n400 ), .A0N(\U1/n489 ), 
        .Y(\U1/n864 ) );
  XOR2_X0P5M_A12TL \U1/U667  ( .A(\U1/key [85]), .B(Din[85]), .Y(\U1/n488 ) );
  AOI22_X0P5M_A12TL \U1/U666  ( .A0(\U1/n1097 ), .A1(\U1/n488 ), .B0(
        \U1/dat_next [85]), .B1(\U1/n404 ), .Y(\U1/n487 ) );
  AO1B2_X0P5M_A12TL \U1/U665  ( .B0(Dout[85]), .B1(\U1/n400 ), .A0N(\U1/n487 ), 
        .Y(\U1/n863 ) );
  XOR2_X0P5M_A12TL \U1/U664  ( .A(\U1/key [86]), .B(Din[86]), .Y(\U1/n486 ) );
  AOI22_X0P5M_A12TL \U1/U663  ( .A0(\U1/n1097 ), .A1(\U1/n486 ), .B0(
        \U1/dat_next [86]), .B1(\U1/n404 ), .Y(\U1/n485 ) );
  AO1B2_X0P5M_A12TL \U1/U662  ( .B0(Dout[86]), .B1(\U1/n400 ), .A0N(\U1/n485 ), 
        .Y(\U1/n862 ) );
  XOR2_X0P5M_A12TL \U1/U661  ( .A(\U1/key [87]), .B(Din[87]), .Y(\U1/n484 ) );
  AOI22_X0P5M_A12TL \U1/U660  ( .A0(\U1/n1097 ), .A1(\U1/n484 ), .B0(
        \U1/dat_next [87]), .B1(\U1/n670 ), .Y(\U1/n483 ) );
  AO1B2_X0P5M_A12TL \U1/U659  ( .B0(Dout[87]), .B1(\U1/n1098 ), .A0N(\U1/n483 ), .Y(\U1/n861 ) );
  XOR2_X0P5M_A12TL \U1/U658  ( .A(\U1/key [88]), .B(Din[88]), .Y(\U1/n482 ) );
  AOI22_X0P5M_A12TL \U1/U657  ( .A0(\U1/n1097 ), .A1(\U1/n482 ), .B0(
        \U1/dat_next [88]), .B1(\U1/n404 ), .Y(\U1/n481 ) );
  AO1B2_X0P5M_A12TL \U1/U656  ( .B0(Dout[88]), .B1(\U1/n1098 ), .A0N(\U1/n481 ), .Y(\U1/n860 ) );
  XOR2_X0P5M_A12TL \U1/U655  ( .A(\U1/key [89]), .B(Din[89]), .Y(\U1/n480 ) );
  AOI22_X0P5M_A12TL \U1/U654  ( .A0(\U1/n1097 ), .A1(\U1/n480 ), .B0(
        \U1/dat_next [89]), .B1(\U1/n404 ), .Y(\U1/n479 ) );
  AO1B2_X0P5M_A12TL \U1/U653  ( .B0(Dout[89]), .B1(\U1/n400 ), .A0N(\U1/n479 ), 
        .Y(\U1/n859 ) );
  XOR2_X0P5M_A12TL \U1/U652  ( .A(\U1/key [90]), .B(Din[90]), .Y(\U1/n478 ) );
  AOI22_X0P5M_A12TL \U1/U651  ( .A0(\U1/n1097 ), .A1(\U1/n478 ), .B0(
        \U1/dat_next [90]), .B1(\U1/n404 ), .Y(\U1/n477 ) );
  AO1B2_X0P5M_A12TL \U1/U650  ( .B0(Dout[90]), .B1(\U1/n400 ), .A0N(\U1/n477 ), 
        .Y(\U1/n858 ) );
  XOR2_X0P5M_A12TL \U1/U649  ( .A(\U1/key [91]), .B(Din[91]), .Y(\U1/n476 ) );
  AOI22_X0P5M_A12TL \U1/U648  ( .A0(\U1/n1097 ), .A1(\U1/n476 ), .B0(
        \U1/dat_next [91]), .B1(\U1/n404 ), .Y(\U1/n475 ) );
  AO1B2_X0P5M_A12TL \U1/U647  ( .B0(Dout[91]), .B1(\U1/n400 ), .A0N(\U1/n475 ), 
        .Y(\U1/n857 ) );
  XOR2_X0P5M_A12TL \U1/U646  ( .A(\U1/key [92]), .B(Din[92]), .Y(\U1/n474 ) );
  AOI22_X0P5M_A12TL \U1/U645  ( .A0(\U1/n1097 ), .A1(\U1/n474 ), .B0(
        \U1/dat_next [92]), .B1(\U1/n404 ), .Y(\U1/n473 ) );
  AO1B2_X0P5M_A12TL \U1/U644  ( .B0(Dout[92]), .B1(\U1/n400 ), .A0N(\U1/n473 ), 
        .Y(\U1/n856 ) );
  XOR2_X0P5M_A12TL \U1/U643  ( .A(\U1/key [93]), .B(Din[93]), .Y(\U1/n472 ) );
  AOI22_X0P5M_A12TL \U1/U642  ( .A0(\U1/n1097 ), .A1(\U1/n472 ), .B0(
        \U1/dat_next [93]), .B1(\U1/n404 ), .Y(\U1/n471 ) );
  AO1B2_X0P5M_A12TL \U1/U641  ( .B0(Dout[93]), .B1(\U1/n400 ), .A0N(\U1/n471 ), 
        .Y(\U1/n855 ) );
  XOR2_X0P5M_A12TL \U1/U640  ( .A(\U1/key [94]), .B(Din[94]), .Y(\U1/n470 ) );
  AOI22_X0P5M_A12TL \U1/U639  ( .A0(\U1/n1097 ), .A1(\U1/n470 ), .B0(
        \U1/dat_next [94]), .B1(\U1/n670 ), .Y(\U1/n469 ) );
  AO1B2_X0P5M_A12TL \U1/U638  ( .B0(Dout[94]), .B1(\U1/n400 ), .A0N(\U1/n469 ), 
        .Y(\U1/n854 ) );
  XOR2_X0P5M_A12TL \U1/U637  ( .A(\U1/key [95]), .B(Din[95]), .Y(\U1/n468 ) );
  AOI22_X0P5M_A12TL \U1/U636  ( .A0(\U1/n1097 ), .A1(\U1/n468 ), .B0(
        \U1/dat_next [95]), .B1(\U1/n404 ), .Y(\U1/n467 ) );
  AO1B2_X0P5M_A12TL \U1/U635  ( .B0(Dout[95]), .B1(\U1/n400 ), .A0N(\U1/n467 ), 
        .Y(\U1/n853 ) );
  XOR2_X0P5M_A12TL \U1/U634  ( .A(\U1/key [96]), .B(Din[96]), .Y(\U1/n466 ) );
  AOI22_X0P5M_A12TL \U1/U633  ( .A0(\U1/n1097 ), .A1(\U1/n466 ), .B0(
        \U1/dat_next [96]), .B1(\U1/n670 ), .Y(\U1/n465 ) );
  AO1B2_X0P5M_A12TL \U1/U632  ( .B0(Dout[96]), .B1(\U1/n400 ), .A0N(\U1/n465 ), 
        .Y(\U1/n852 ) );
  XOR2_X0P5M_A12TL \U1/U631  ( .A(\U1/key [97]), .B(Din[97]), .Y(\U1/n464 ) );
  AOI22_X0P5M_A12TL \U1/U630  ( .A0(\U1/n1097 ), .A1(\U1/n464 ), .B0(
        \U1/dat_next [97]), .B1(\U1/n670 ), .Y(\U1/n463 ) );
  AO1B2_X0P5M_A12TL \U1/U629  ( .B0(Dout[97]), .B1(\U1/n400 ), .A0N(\U1/n463 ), 
        .Y(\U1/n851 ) );
  XOR2_X0P5M_A12TL \U1/U628  ( .A(\U1/key [98]), .B(Din[98]), .Y(\U1/n462 ) );
  AOI22_X0P5M_A12TL \U1/U627  ( .A0(\U1/n1097 ), .A1(\U1/n462 ), .B0(
        \U1/dat_next [98]), .B1(\U1/n670 ), .Y(\U1/n461 ) );
  AO1B2_X0P5M_A12TL \U1/U626  ( .B0(Dout[98]), .B1(\U1/n400 ), .A0N(\U1/n461 ), 
        .Y(\U1/n850 ) );
  XOR2_X0P5M_A12TL \U1/U625  ( .A(\U1/key [99]), .B(Din[99]), .Y(\U1/n460 ) );
  AOI22_X0P5M_A12TL \U1/U624  ( .A0(\U1/n1097 ), .A1(\U1/n460 ), .B0(
        \U1/dat_next [99]), .B1(\U1/n670 ), .Y(\U1/n459 ) );
  AO1B2_X0P5M_A12TL \U1/U623  ( .B0(Dout[99]), .B1(\U1/n400 ), .A0N(\U1/n459 ), 
        .Y(\U1/n849 ) );
  XOR2_X0P5M_A12TL \U1/U622  ( .A(\U1/key [100]), .B(Din[100]), .Y(\U1/n458 )
         );
  AOI22_X0P5M_A12TL \U1/U621  ( .A0(\U1/n1097 ), .A1(\U1/n458 ), .B0(
        \U1/dat_next [100]), .B1(\U1/n404 ), .Y(\U1/n457 ) );
  AO1B2_X0P5M_A12TL \U1/U620  ( .B0(Dout[100]), .B1(\U1/n400 ), .A0N(\U1/n457 ), .Y(\U1/n848 ) );
  XOR2_X0P5M_A12TL \U1/U619  ( .A(\U1/key [101]), .B(Din[101]), .Y(\U1/n456 )
         );
  AOI22_X0P5M_A12TL \U1/U618  ( .A0(\U1/n1097 ), .A1(\U1/n456 ), .B0(
        \U1/dat_next [101]), .B1(\U1/n670 ), .Y(\U1/n455 ) );
  AO1B2_X0P5M_A12TL \U1/U617  ( .B0(Dout[101]), .B1(\U1/n400 ), .A0N(\U1/n455 ), .Y(\U1/n847 ) );
  XOR2_X0P5M_A12TL \U1/U616  ( .A(\U1/key [102]), .B(Din[102]), .Y(\U1/n454 )
         );
  AOI22_X0P5M_A12TL \U1/U615  ( .A0(\U1/n1097 ), .A1(\U1/n454 ), .B0(
        \U1/dat_next [102]), .B1(\U1/n404 ), .Y(\U1/n453 ) );
  AO1B2_X0P5M_A12TL \U1/U614  ( .B0(Dout[102]), .B1(\U1/n400 ), .A0N(\U1/n453 ), .Y(\U1/n846 ) );
  XOR2_X0P5M_A12TL \U1/U613  ( .A(\U1/key [103]), .B(Din[103]), .Y(\U1/n452 )
         );
  AOI22_X0P5M_A12TL \U1/U612  ( .A0(\U1/n1097 ), .A1(\U1/n452 ), .B0(
        \U1/dat_next [103]), .B1(\U1/n670 ), .Y(\U1/n451 ) );
  AO1B2_X0P5M_A12TL \U1/U611  ( .B0(Dout[103]), .B1(\U1/n1098 ), .A0N(
        \U1/n451 ), .Y(\U1/n845 ) );
  XOR2_X0P5M_A12TL \U1/U610  ( .A(\U1/key [104]), .B(Din[104]), .Y(\U1/n450 )
         );
  AOI22_X0P5M_A12TL \U1/U609  ( .A0(\U1/n402 ), .A1(\U1/n450 ), .B0(
        \U1/dat_next [104]), .B1(\U1/n670 ), .Y(\U1/n449 ) );
  AO1B2_X0P5M_A12TL \U1/U608  ( .B0(Dout[104]), .B1(\U1/n1098 ), .A0N(
        \U1/n449 ), .Y(\U1/n844 ) );
  XOR2_X0P5M_A12TL \U1/U607  ( .A(\U1/key [105]), .B(Din[105]), .Y(\U1/n448 )
         );
  AOI22_X0P5M_A12TL \U1/U606  ( .A0(\U1/n402 ), .A1(\U1/n448 ), .B0(
        \U1/dat_next [105]), .B1(\U1/n670 ), .Y(\U1/n447 ) );
  AO1B2_X0P5M_A12TL \U1/U605  ( .B0(Dout[105]), .B1(\U1/n400 ), .A0N(\U1/n447 ), .Y(\U1/n843 ) );
  XOR2_X0P5M_A12TL \U1/U604  ( .A(\U1/key [106]), .B(Din[106]), .Y(\U1/n446 )
         );
  AOI22_X0P5M_A12TL \U1/U603  ( .A0(\U1/n402 ), .A1(\U1/n446 ), .B0(
        \U1/dat_next [106]), .B1(\U1/n670 ), .Y(\U1/n445 ) );
  AO1B2_X0P5M_A12TL \U1/U602  ( .B0(Dout[106]), .B1(\U1/n400 ), .A0N(\U1/n445 ), .Y(\U1/n842 ) );
  XOR2_X0P5M_A12TL \U1/U601  ( .A(\U1/key [107]), .B(Din[107]), .Y(\U1/n444 )
         );
  AOI22_X0P5M_A12TL \U1/U600  ( .A0(\U1/n402 ), .A1(\U1/n444 ), .B0(
        \U1/dat_next [107]), .B1(\U1/n670 ), .Y(\U1/n443 ) );
  AO1B2_X0P5M_A12TL \U1/U599  ( .B0(Dout[107]), .B1(\U1/n400 ), .A0N(\U1/n443 ), .Y(\U1/n841 ) );
  XOR2_X0P5M_A12TL \U1/U598  ( .A(\U1/key [108]), .B(Din[108]), .Y(\U1/n442 )
         );
  AOI22_X0P5M_A12TL \U1/U597  ( .A0(\U1/n402 ), .A1(\U1/n442 ), .B0(
        \U1/dat_next [108]), .B1(\U1/n670 ), .Y(\U1/n441 ) );
  AO1B2_X0P5M_A12TL \U1/U596  ( .B0(Dout[108]), .B1(\U1/n400 ), .A0N(\U1/n441 ), .Y(\U1/n840 ) );
  XOR2_X0P5M_A12TL \U1/U595  ( .A(\U1/key [109]), .B(Din[109]), .Y(\U1/n440 )
         );
  AOI22_X0P5M_A12TL \U1/U594  ( .A0(\U1/n402 ), .A1(\U1/n440 ), .B0(
        \U1/dat_next [109]), .B1(\U1/n670 ), .Y(\U1/n439 ) );
  AO1B2_X0P5M_A12TL \U1/U593  ( .B0(Dout[109]), .B1(\U1/n400 ), .A0N(\U1/n439 ), .Y(\U1/n839 ) );
  XOR2_X0P5M_A12TL \U1/U592  ( .A(\U1/key [110]), .B(Din[110]), .Y(\U1/n438 )
         );
  AOI22_X0P5M_A12TL \U1/U591  ( .A0(\U1/n402 ), .A1(\U1/n438 ), .B0(
        \U1/dat_next [110]), .B1(\U1/n670 ), .Y(\U1/n437 ) );
  AO1B2_X0P5M_A12TL \U1/U590  ( .B0(Dout[110]), .B1(\U1/n400 ), .A0N(\U1/n437 ), .Y(\U1/n838 ) );
  XOR2_X0P5M_A12TL \U1/U589  ( .A(\U1/key [111]), .B(Din[111]), .Y(\U1/n436 )
         );
  AOI22_X0P5M_A12TL \U1/U588  ( .A0(\U1/n402 ), .A1(\U1/n436 ), .B0(
        \U1/dat_next [111]), .B1(\U1/n670 ), .Y(\U1/n435 ) );
  AO1B2_X0P5M_A12TL \U1/U587  ( .B0(Dout[111]), .B1(\U1/n400 ), .A0N(\U1/n435 ), .Y(\U1/n837 ) );
  XOR2_X0P5M_A12TL \U1/U586  ( .A(\U1/key [112]), .B(Din[112]), .Y(\U1/n434 )
         );
  AOI22_X0P5M_A12TL \U1/U585  ( .A0(\U1/n1097 ), .A1(\U1/n434 ), .B0(
        \U1/dat_next [112]), .B1(\U1/n404 ), .Y(\U1/n433 ) );
  AO1B2_X0P5M_A12TL \U1/U584  ( .B0(Dout[112]), .B1(\U1/n400 ), .A0N(\U1/n433 ), .Y(\U1/n836 ) );
  XOR2_X0P5M_A12TL \U1/U583  ( .A(\U1/key [113]), .B(Din[113]), .Y(\U1/n432 )
         );
  AOI22_X0P5M_A12TL \U1/U582  ( .A0(\U1/n1097 ), .A1(\U1/n432 ), .B0(
        \U1/dat_next [113]), .B1(\U1/n670 ), .Y(\U1/n431 ) );
  AO1B2_X0P5M_A12TL \U1/U581  ( .B0(Dout[113]), .B1(\U1/n400 ), .A0N(\U1/n431 ), .Y(\U1/n835 ) );
  XOR2_X0P5M_A12TL \U1/U580  ( .A(\U1/key [114]), .B(Din[114]), .Y(\U1/n430 )
         );
  AOI22_X0P5M_A12TL \U1/U579  ( .A0(\U1/n1097 ), .A1(\U1/n430 ), .B0(
        \U1/dat_next [114]), .B1(\U1/n670 ), .Y(\U1/n429 ) );
  AO1B2_X0P5M_A12TL \U1/U578  ( .B0(Dout[114]), .B1(\U1/n400 ), .A0N(\U1/n429 ), .Y(\U1/n834 ) );
  XOR2_X0P5M_A12TL \U1/U577  ( .A(\U1/key [115]), .B(Din[115]), .Y(\U1/n428 )
         );
  AOI22_X0P5M_A12TL \U1/U576  ( .A0(\U1/n1097 ), .A1(\U1/n428 ), .B0(
        \U1/dat_next [115]), .B1(\U1/n404 ), .Y(\U1/n427 ) );
  AO1B2_X0P5M_A12TL \U1/U575  ( .B0(Dout[115]), .B1(\U1/n400 ), .A0N(\U1/n427 ), .Y(\U1/n833 ) );
  XOR2_X0P5M_A12TL \U1/U574  ( .A(\U1/key [116]), .B(Din[116]), .Y(\U1/n426 )
         );
  AOI22_X0P5M_A12TL \U1/U573  ( .A0(\U1/n1097 ), .A1(\U1/n426 ), .B0(
        \U1/dat_next [116]), .B1(\U1/n404 ), .Y(\U1/n425 ) );
  AO1B2_X0P5M_A12TL \U1/U572  ( .B0(Dout[116]), .B1(\U1/n400 ), .A0N(\U1/n425 ), .Y(\U1/n832 ) );
  XOR2_X0P5M_A12TL \U1/U571  ( .A(\U1/key [117]), .B(Din[117]), .Y(\U1/n424 )
         );
  AOI22_X0P5M_A12TL \U1/U570  ( .A0(\U1/n1097 ), .A1(\U1/n424 ), .B0(
        \U1/dat_next [117]), .B1(\U1/n404 ), .Y(\U1/n423 ) );
  AO1B2_X0P5M_A12TL \U1/U569  ( .B0(Dout[117]), .B1(\U1/n400 ), .A0N(\U1/n423 ), .Y(\U1/n831 ) );
  XOR2_X0P5M_A12TL \U1/U568  ( .A(\U1/key [118]), .B(Din[118]), .Y(\U1/n422 )
         );
  AOI22_X0P5M_A12TL \U1/U567  ( .A0(\U1/n1097 ), .A1(\U1/n422 ), .B0(
        \U1/dat_next [118]), .B1(\U1/n404 ), .Y(\U1/n421 ) );
  AO1B2_X0P5M_A12TL \U1/U566  ( .B0(Dout[118]), .B1(\U1/n400 ), .A0N(\U1/n421 ), .Y(\U1/n830 ) );
  XOR2_X0P5M_A12TL \U1/U565  ( .A(\U1/key [119]), .B(Din[119]), .Y(\U1/n420 )
         );
  AOI22_X0P5M_A12TL \U1/U564  ( .A0(\U1/n1097 ), .A1(\U1/n420 ), .B0(
        \U1/dat_next [119]), .B1(\U1/n404 ), .Y(\U1/n419 ) );
  AO1B2_X0P5M_A12TL \U1/U563  ( .B0(Dout[119]), .B1(\U1/n400 ), .A0N(\U1/n419 ), .Y(\U1/n829 ) );
  XOR2_X0P5M_A12TL \U1/U562  ( .A(\U1/key [120]), .B(Din[120]), .Y(\U1/n418 )
         );
  AOI22_X0P5M_A12TL \U1/U561  ( .A0(\U1/n1097 ), .A1(\U1/n418 ), .B0(
        \U1/dat_next [120]), .B1(\U1/n404 ), .Y(\U1/n417 ) );
  AO1B2_X0P5M_A12TL \U1/U560  ( .B0(Dout[120]), .B1(\U1/n400 ), .A0N(\U1/n417 ), .Y(\U1/n828 ) );
  XOR2_X0P5M_A12TL \U1/U559  ( .A(\U1/key [121]), .B(Din[121]), .Y(\U1/n416 )
         );
  AOI22_X0P5M_A12TL \U1/U558  ( .A0(\U1/n1097 ), .A1(\U1/n416 ), .B0(
        \U1/dat_next [121]), .B1(\U1/n404 ), .Y(\U1/n415 ) );
  AO1B2_X0P5M_A12TL \U1/U557  ( .B0(Dout[121]), .B1(\U1/n400 ), .A0N(\U1/n415 ), .Y(\U1/n827 ) );
  XOR2_X0P5M_A12TL \U1/U556  ( .A(\U1/key [122]), .B(Din[122]), .Y(\U1/n414 )
         );
  AOI22_X0P5M_A12TL \U1/U555  ( .A0(\U1/n1097 ), .A1(\U1/n414 ), .B0(
        \U1/dat_next [122]), .B1(\U1/n404 ), .Y(\U1/n413 ) );
  AO1B2_X0P5M_A12TL \U1/U554  ( .B0(Dout[122]), .B1(\U1/n400 ), .A0N(\U1/n413 ), .Y(\U1/n826 ) );
  XOR2_X0P5M_A12TL \U1/U553  ( .A(\U1/key [123]), .B(Din[123]), .Y(\U1/n412 )
         );
  AOI22_X0P5M_A12TL \U1/U552  ( .A0(\U1/n1097 ), .A1(\U1/n412 ), .B0(
        \U1/dat_next [123]), .B1(\U1/n404 ), .Y(\U1/n411 ) );
  AO1B2_X0P5M_A12TL \U1/U551  ( .B0(Dout[123]), .B1(\U1/n400 ), .A0N(\U1/n411 ), .Y(\U1/n825 ) );
  XOR2_X0P5M_A12TL \U1/U550  ( .A(\U1/key [124]), .B(Din[124]), .Y(\U1/n410 )
         );
  AOI22_X0P5M_A12TL \U1/U549  ( .A0(\U1/n1097 ), .A1(\U1/n410 ), .B0(
        \U1/dat_next [124]), .B1(\U1/n404 ), .Y(\U1/n409 ) );
  AO1B2_X0P5M_A12TL \U1/U548  ( .B0(Dout[124]), .B1(\U1/n400 ), .A0N(\U1/n409 ), .Y(\U1/n824 ) );
  XOR2_X0P5M_A12TL \U1/U547  ( .A(\U1/key [125]), .B(Din[125]), .Y(\U1/n408 )
         );
  AOI22_X0P5M_A12TL \U1/U546  ( .A0(\U1/n1097 ), .A1(\U1/n408 ), .B0(
        \U1/dat_next [125]), .B1(\U1/n404 ), .Y(\U1/n407 ) );
  AO1B2_X0P5M_A12TL \U1/U545  ( .B0(Dout[125]), .B1(\U1/n1098 ), .A0N(
        \U1/n407 ), .Y(\U1/n823 ) );
  XOR2_X0P5M_A12TL \U1/U544  ( .A(\U1/key [126]), .B(Din[126]), .Y(\U1/n406 )
         );
  AOI22_X0P5M_A12TL \U1/U543  ( .A0(\U1/n1097 ), .A1(\U1/n406 ), .B0(
        \U1/dat_next [126]), .B1(\U1/n404 ), .Y(\U1/n405 ) );
  AO1B2_X0P5M_A12TL \U1/U542  ( .B0(Dout[126]), .B1(\U1/n1098 ), .A0N(
        \U1/n405 ), .Y(\U1/n822 ) );
  XOR2_X0P5M_A12TL \U1/U541  ( .A(\U1/key [127]), .B(Din[127]), .Y(\U1/n403 )
         );
  AOI22_X0P5M_A12TL \U1/U540  ( .A0(\U1/n1097 ), .A1(\U1/n403 ), .B0(
        \U1/dat_next [127]), .B1(\U1/n404 ), .Y(\U1/n401 ) );
  AO1B2_X0P5M_A12TL \U1/U539  ( .B0(Dout[127]), .B1(\U1/n1098 ), .A0N(
        \U1/n401 ), .Y(\U1/n821 ) );
  OAI2XB1_X0P5M_A12TL \U1/U538  ( .A1N(Kvld), .A0(EN), .B0(\U1/n1105 ), .Y(
        \U1/n820 ) );
  AO22_X0P5M_A12TL \U1/U537  ( .A0(EN), .A1(\U1/rnd [9]), .B0(\U1/n1099 ), 
        .B1(\U1/sel ), .Y(\U1/n811 ) );
  AO22_X0P5M_A12TL \U1/U536  ( .A0(\U1/sel ), .A1(EN), .B0(Dvld), .B1(
        \U1/n1099 ), .Y(\U1/n810 ) );
  INV_X0P5B_A12TL \U1/U535  ( .A(\U1/n819 ), .Y(\U1/n398 ) );
  INV_X0P5B_A12TL \U1/U534  ( .A(\U1/n818 ), .Y(\U1/n399 ) );
  OR6_X0P5M_A12TL \U1/U533  ( .A(\U1/n1099 ), .B(\U1/n398 ), .C(\U1/n399 ), 
        .D(\U1/sel ), .E(\U1/rnd [9]), .F(KDrdy2), .Y(\U1/n390 ) );
  INV_X0P5B_A12TL \U1/U532  ( .A(\U1/n814 ), .Y(\U1/n392 ) );
  INV_X0P5B_A12TL \U1/U531  ( .A(\U1/n813 ), .Y(\U1/n393 ) );
  INV_X0P5B_A12TL \U1/U530  ( .A(\U1/n812 ), .Y(\U1/n394 ) );
  INV_X0P5B_A12TL \U1/U529  ( .A(\U1/n817 ), .Y(\U1/n395 ) );
  INV_X0P5B_A12TL \U1/U528  ( .A(\U1/n816 ), .Y(\U1/n396 ) );
  INV_X0P5B_A12TL \U1/U527  ( .A(\U1/n815 ), .Y(\U1/n397 ) );
  OR6_X0P5M_A12TL \U1/U526  ( .A(\U1/n392 ), .B(\U1/n393 ), .C(\U1/n394 ), .D(
        \U1/n395 ), .E(\U1/n396 ), .F(\U1/n397 ), .Y(\U1/n391 ) );
  OA22_X0P5M_A12TL \U1/U525  ( .A0(\U1/n390 ), .A1(\U1/n391 ), .B0(EN), .B1(
        BSY), .Y(\U1/n809 ) );
  INV_X0P5B_A12TL \U1/U524  ( .A(Kin[0]), .Y(\U1/n386 ) );
  NAND2_X0P5A_A12TL \U1/U523  ( .A(\U1/rkey [0]), .B(\U1/n7 ), .Y(\U1/n387 )
         );
  NOR3_X0P5A_A12TL \U1/U522  ( .A(\U1/n1099 ), .B(KDrdy), .C(\U1/n389 ), .Y(
        \U1/n5 ) );
  NOR3_X0P5A_A12TL \U1/U521  ( .A(KDrdy), .B(\U1/rnd [0]), .C(\U1/n7 ), .Y(
        \U1/n6 ) );
  AOI22_X0P5M_A12TL \U1/U520  ( .A0(\U1/key [0]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [0]), .B1(\U1/n1101 ), .Y(\U1/n388 ) );
  OAI211_X0P5M_A12TL \U1/U519  ( .A0(\U1/n1106 ), .A1(\U1/n386 ), .B0(
        \U1/n387 ), .C0(\U1/n388 ), .Y(\U1/n801 ) );
  INV_X0P5B_A12TL \U1/U518  ( .A(Kin[1]), .Y(\U1/n383 ) );
  NAND2_X0P5A_A12TL \U1/U517  ( .A(\U1/rkey [1]), .B(\U1/n7 ), .Y(\U1/n384 )
         );
  AOI22_X0P5M_A12TL \U1/U516  ( .A0(\U1/key [1]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [1]), .B1(\U1/n1101 ), .Y(\U1/n385 ) );
  OAI211_X0P5M_A12TL \U1/U515  ( .A0(\U1/n1107 ), .A1(\U1/n383 ), .B0(
        \U1/n384 ), .C0(\U1/n385 ), .Y(\U1/n800 ) );
  INV_X0P5B_A12TL \U1/U514  ( .A(Kin[2]), .Y(\U1/n380 ) );
  NAND2_X0P5A_A12TL \U1/U513  ( .A(\U1/rkey [2]), .B(\U1/n7 ), .Y(\U1/n381 )
         );
  AOI22_X0P5M_A12TL \U1/U512  ( .A0(\U1/key [2]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [2]), .B1(\U1/n1101 ), .Y(\U1/n382 ) );
  OAI211_X0P5M_A12TL \U1/U511  ( .A0(\U1/n1106 ), .A1(\U1/n380 ), .B0(
        \U1/n381 ), .C0(\U1/n382 ), .Y(\U1/n799 ) );
  INV_X0P5B_A12TL \U1/U510  ( .A(Kin[3]), .Y(\U1/n377 ) );
  NAND2_X0P5A_A12TL \U1/U509  ( .A(\U1/rkey [3]), .B(\U1/n7 ), .Y(\U1/n378 )
         );
  AOI22_X0P5M_A12TL \U1/U508  ( .A0(\U1/key [3]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [3]), .B1(\U1/n1101 ), .Y(\U1/n379 ) );
  OAI211_X0P5M_A12TL \U1/U507  ( .A0(\U1/n1107 ), .A1(\U1/n377 ), .B0(
        \U1/n378 ), .C0(\U1/n379 ), .Y(\U1/n798 ) );
  INV_X0P5B_A12TL \U1/U506  ( .A(Kin[4]), .Y(\U1/n374 ) );
  NAND2_X0P5A_A12TL \U1/U505  ( .A(\U1/rkey [4]), .B(\U1/n7 ), .Y(\U1/n375 )
         );
  AOI22_X0P5M_A12TL \U1/U504  ( .A0(\U1/key [4]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [4]), .B1(\U1/n1101 ), .Y(\U1/n376 ) );
  OAI211_X0P5M_A12TL \U1/U503  ( .A0(\U1/n1105 ), .A1(\U1/n374 ), .B0(
        \U1/n375 ), .C0(\U1/n376 ), .Y(\U1/n797 ) );
  INV_X0P5B_A12TL \U1/U502  ( .A(Kin[5]), .Y(\U1/n371 ) );
  NAND2_X0P5A_A12TL \U1/U501  ( .A(\U1/rkey [5]), .B(\U1/n7 ), .Y(\U1/n372 )
         );
  AOI22_X0P5M_A12TL \U1/U500  ( .A0(\U1/key [5]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [5]), .B1(\U1/n1101 ), .Y(\U1/n373 ) );
  OAI211_X0P5M_A12TL \U1/U499  ( .A0(\U1/n1106 ), .A1(\U1/n371 ), .B0(
        \U1/n372 ), .C0(\U1/n373 ), .Y(\U1/n796 ) );
  INV_X0P5B_A12TL \U1/U498  ( .A(Kin[6]), .Y(\U1/n368 ) );
  NAND2_X0P5A_A12TL \U1/U497  ( .A(\U1/rkey [6]), .B(\U1/n1099 ), .Y(\U1/n369 ) );
  AOI22_X0P5M_A12TL \U1/U496  ( .A0(\U1/key [6]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [6]), .B1(\U1/n1101 ), .Y(\U1/n370 ) );
  OAI211_X0P5M_A12TL \U1/U495  ( .A0(\U1/n1107 ), .A1(\U1/n368 ), .B0(
        \U1/n369 ), .C0(\U1/n370 ), .Y(\U1/n795 ) );
  INV_X0P5B_A12TL \U1/U494  ( .A(Kin[7]), .Y(\U1/n365 ) );
  NAND2_X0P5A_A12TL \U1/U493  ( .A(\U1/rkey [7]), .B(\U1/n1099 ), .Y(\U1/n366 ) );
  AOI22_X0P5M_A12TL \U1/U492  ( .A0(\U1/key [7]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [7]), .B1(\U1/n1101 ), .Y(\U1/n367 ) );
  OAI211_X0P5M_A12TL \U1/U491  ( .A0(\U1/n1107 ), .A1(\U1/n365 ), .B0(
        \U1/n366 ), .C0(\U1/n367 ), .Y(\U1/n794 ) );
  INV_X0P5B_A12TL \U1/U490  ( .A(Kin[8]), .Y(\U1/n362 ) );
  NAND2_X0P5A_A12TL \U1/U489  ( .A(\U1/rkey [8]), .B(\U1/n1099 ), .Y(\U1/n363 ) );
  AOI22_X0P5M_A12TL \U1/U488  ( .A0(\U1/key [8]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [8]), .B1(\U1/n1101 ), .Y(\U1/n364 ) );
  OAI211_X0P5M_A12TL \U1/U487  ( .A0(\U1/n1107 ), .A1(\U1/n362 ), .B0(
        \U1/n363 ), .C0(\U1/n364 ), .Y(\U1/n793 ) );
  INV_X0P5B_A12TL \U1/U486  ( .A(Kin[9]), .Y(\U1/n359 ) );
  NAND2_X0P5A_A12TL \U1/U485  ( .A(\U1/rkey [9]), .B(\U1/n1099 ), .Y(\U1/n360 ) );
  AOI22_X0P5M_A12TL \U1/U484  ( .A0(\U1/key [9]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [9]), .B1(\U1/n1101 ), .Y(\U1/n361 ) );
  OAI211_X0P5M_A12TL \U1/U483  ( .A0(\U1/n1107 ), .A1(\U1/n359 ), .B0(
        \U1/n360 ), .C0(\U1/n361 ), .Y(\U1/n792 ) );
  INV_X0P5B_A12TL \U1/U482  ( .A(Kin[10]), .Y(\U1/n356 ) );
  NAND2_X0P5A_A12TL \U1/U481  ( .A(\U1/rkey [10]), .B(\U1/n1099 ), .Y(
        \U1/n357 ) );
  AOI22_X0P5M_A12TL \U1/U480  ( .A0(\U1/key [10]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [10]), .B1(\U1/n1100 ), .Y(\U1/n358 ) );
  OAI211_X0P5M_A12TL \U1/U479  ( .A0(\U1/n1107 ), .A1(\U1/n356 ), .B0(
        \U1/n357 ), .C0(\U1/n358 ), .Y(\U1/n791 ) );
  INV_X0P5B_A12TL \U1/U478  ( .A(Kin[11]), .Y(\U1/n353 ) );
  NAND2_X0P5A_A12TL \U1/U477  ( .A(\U1/rkey [11]), .B(\U1/n1099 ), .Y(
        \U1/n354 ) );
  AOI22_X0P5M_A12TL \U1/U476  ( .A0(\U1/key [11]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [11]), .B1(\U1/n1101 ), .Y(\U1/n355 ) );
  OAI211_X0P5M_A12TL \U1/U475  ( .A0(\U1/n1107 ), .A1(\U1/n353 ), .B0(
        \U1/n354 ), .C0(\U1/n355 ), .Y(\U1/n790 ) );
  INV_X0P5B_A12TL \U1/U474  ( .A(Kin[12]), .Y(\U1/n350 ) );
  NAND2_X0P5A_A12TL \U1/U473  ( .A(\U1/rkey [12]), .B(\U1/n7 ), .Y(\U1/n351 )
         );
  AOI22_X0P5M_A12TL \U1/U472  ( .A0(\U1/key [12]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [12]), .B1(\U1/n1101 ), .Y(\U1/n352 ) );
  OAI211_X0P5M_A12TL \U1/U471  ( .A0(\U1/n1107 ), .A1(\U1/n350 ), .B0(
        \U1/n351 ), .C0(\U1/n352 ), .Y(\U1/n789 ) );
  INV_X0P5B_A12TL \U1/U470  ( .A(Kin[13]), .Y(\U1/n347 ) );
  NAND2_X0P5A_A12TL \U1/U469  ( .A(\U1/rkey [13]), .B(\U1/n7 ), .Y(\U1/n348 )
         );
  AOI22_X0P5M_A12TL \U1/U468  ( .A0(\U1/key [13]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [13]), .B1(\U1/n1101 ), .Y(\U1/n349 ) );
  OAI211_X0P5M_A12TL \U1/U467  ( .A0(\U1/n1107 ), .A1(\U1/n347 ), .B0(
        \U1/n348 ), .C0(\U1/n349 ), .Y(\U1/n788 ) );
  INV_X0P5B_A12TL \U1/U466  ( .A(Kin[14]), .Y(\U1/n344 ) );
  NAND2_X0P5A_A12TL \U1/U465  ( .A(\U1/rkey [14]), .B(\U1/n7 ), .Y(\U1/n345 )
         );
  AOI22_X0P5M_A12TL \U1/U464  ( .A0(\U1/key [14]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [14]), .B1(\U1/n1101 ), .Y(\U1/n346 ) );
  OAI211_X0P5M_A12TL \U1/U463  ( .A0(\U1/n1107 ), .A1(\U1/n344 ), .B0(
        \U1/n345 ), .C0(\U1/n346 ), .Y(\U1/n787 ) );
  INV_X0P5B_A12TL \U1/U462  ( .A(Kin[15]), .Y(\U1/n341 ) );
  NAND2_X0P5A_A12TL \U1/U461  ( .A(\U1/rkey [15]), .B(\U1/n7 ), .Y(\U1/n342 )
         );
  AOI22_X0P5M_A12TL \U1/U460  ( .A0(\U1/key [15]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [15]), .B1(\U1/n1101 ), .Y(\U1/n343 ) );
  OAI211_X0P5M_A12TL \U1/U459  ( .A0(\U1/n1107 ), .A1(\U1/n341 ), .B0(
        \U1/n342 ), .C0(\U1/n343 ), .Y(\U1/n786 ) );
  INV_X0P5B_A12TL \U1/U458  ( .A(Kin[16]), .Y(\U1/n338 ) );
  NAND2_X0P5A_A12TL \U1/U457  ( .A(\U1/rkey [16]), .B(\U1/n1099 ), .Y(
        \U1/n339 ) );
  AOI22_X0P5M_A12TL \U1/U456  ( .A0(\U1/key [16]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [16]), .B1(\U1/n1101 ), .Y(\U1/n340 ) );
  OAI211_X0P5M_A12TL \U1/U455  ( .A0(\U1/n1107 ), .A1(\U1/n338 ), .B0(
        \U1/n339 ), .C0(\U1/n340 ), .Y(\U1/n785 ) );
  INV_X0P5B_A12TL \U1/U454  ( .A(Kin[17]), .Y(\U1/n335 ) );
  NAND2_X0P5A_A12TL \U1/U453  ( .A(\U1/rkey [17]), .B(\U1/n7 ), .Y(\U1/n336 )
         );
  AOI22_X0P5M_A12TL \U1/U452  ( .A0(\U1/key [17]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [17]), .B1(\U1/n1101 ), .Y(\U1/n337 ) );
  OAI211_X0P5M_A12TL \U1/U451  ( .A0(\U1/n1107 ), .A1(\U1/n335 ), .B0(
        \U1/n336 ), .C0(\U1/n337 ), .Y(\U1/n784 ) );
  INV_X0P5B_A12TL \U1/U450  ( .A(Kin[18]), .Y(\U1/n332 ) );
  NAND2_X0P5A_A12TL \U1/U449  ( .A(\U1/rkey [18]), .B(\U1/n1099 ), .Y(
        \U1/n333 ) );
  AOI22_X0P5M_A12TL \U1/U448  ( .A0(\U1/key [18]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [18]), .B1(\U1/n1101 ), .Y(\U1/n334 ) );
  OAI211_X0P5M_A12TL \U1/U447  ( .A0(\U1/n1107 ), .A1(\U1/n332 ), .B0(
        \U1/n333 ), .C0(\U1/n334 ), .Y(\U1/n783 ) );
  INV_X0P5B_A12TL \U1/U446  ( .A(Kin[19]), .Y(\U1/n329 ) );
  NAND2_X0P5A_A12TL \U1/U445  ( .A(\U1/rkey [19]), .B(\U1/n7 ), .Y(\U1/n330 )
         );
  AOI22_X0P5M_A12TL \U1/U444  ( .A0(\U1/key [19]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [19]), .B1(\U1/n1101 ), .Y(\U1/n331 ) );
  OAI211_X0P5M_A12TL \U1/U443  ( .A0(\U1/n1106 ), .A1(\U1/n329 ), .B0(
        \U1/n330 ), .C0(\U1/n331 ), .Y(\U1/n782 ) );
  INV_X0P5B_A12TL \U1/U442  ( .A(Kin[20]), .Y(\U1/n326 ) );
  NAND2_X0P5A_A12TL \U1/U441  ( .A(\U1/rkey [20]), .B(\U1/n7 ), .Y(\U1/n327 )
         );
  AOI22_X0P5M_A12TL \U1/U440  ( .A0(\U1/key [20]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [20]), .B1(\U1/n1101 ), .Y(\U1/n328 ) );
  OAI211_X0P5M_A12TL \U1/U439  ( .A0(\U1/n1106 ), .A1(\U1/n326 ), .B0(
        \U1/n327 ), .C0(\U1/n328 ), .Y(\U1/n781 ) );
  INV_X0P5B_A12TL \U1/U438  ( .A(Kin[21]), .Y(\U1/n323 ) );
  NAND2_X0P5A_A12TL \U1/U437  ( .A(\U1/rkey [21]), .B(\U1/n7 ), .Y(\U1/n324 )
         );
  AOI22_X0P5M_A12TL \U1/U436  ( .A0(\U1/key [21]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [21]), .B1(\U1/n1101 ), .Y(\U1/n325 ) );
  OAI211_X0P5M_A12TL \U1/U435  ( .A0(\U1/n1106 ), .A1(\U1/n323 ), .B0(
        \U1/n324 ), .C0(\U1/n325 ), .Y(\U1/n780 ) );
  INV_X0P5B_A12TL \U1/U434  ( .A(Kin[22]), .Y(\U1/n320 ) );
  NAND2_X0P5A_A12TL \U1/U433  ( .A(\U1/rkey [22]), .B(\U1/n7 ), .Y(\U1/n321 )
         );
  AOI22_X0P5M_A12TL \U1/U432  ( .A0(\U1/key [22]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [22]), .B1(\U1/n1101 ), .Y(\U1/n322 ) );
  OAI211_X0P5M_A12TL \U1/U431  ( .A0(\U1/n1106 ), .A1(\U1/n320 ), .B0(
        \U1/n321 ), .C0(\U1/n322 ), .Y(\U1/n779 ) );
  INV_X0P5B_A12TL \U1/U430  ( .A(Kin[23]), .Y(\U1/n317 ) );
  NAND2_X0P5A_A12TL \U1/U429  ( .A(\U1/rkey [23]), .B(\U1/n7 ), .Y(\U1/n318 )
         );
  AOI22_X0P5M_A12TL \U1/U428  ( .A0(\U1/key [23]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [23]), .B1(\U1/n1101 ), .Y(\U1/n319 ) );
  OAI211_X0P5M_A12TL \U1/U427  ( .A0(\U1/n1106 ), .A1(\U1/n317 ), .B0(
        \U1/n318 ), .C0(\U1/n319 ), .Y(\U1/n778 ) );
  INV_X0P5B_A12TL \U1/U426  ( .A(Kin[24]), .Y(\U1/n314 ) );
  NAND2_X0P5A_A12TL \U1/U425  ( .A(\U1/rkey [24]), .B(\U1/n7 ), .Y(\U1/n315 )
         );
  AOI22_X0P5M_A12TL \U1/U424  ( .A0(\U1/key [24]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [24]), .B1(\U1/n1101 ), .Y(\U1/n316 ) );
  OAI211_X0P5M_A12TL \U1/U423  ( .A0(\U1/n1106 ), .A1(\U1/n314 ), .B0(
        \U1/n315 ), .C0(\U1/n316 ), .Y(\U1/n777 ) );
  INV_X0P5B_A12TL \U1/U422  ( .A(Kin[25]), .Y(\U1/n311 ) );
  NAND2_X0P5A_A12TL \U1/U421  ( .A(\U1/rkey [25]), .B(\U1/n7 ), .Y(\U1/n312 )
         );
  AOI22_X0P5M_A12TL \U1/U420  ( .A0(\U1/key [25]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [25]), .B1(\U1/n1101 ), .Y(\U1/n313 ) );
  OAI211_X0P5M_A12TL \U1/U419  ( .A0(\U1/n1106 ), .A1(\U1/n311 ), .B0(
        \U1/n312 ), .C0(\U1/n313 ), .Y(\U1/n776 ) );
  INV_X0P5B_A12TL \U1/U418  ( .A(Kin[26]), .Y(\U1/n308 ) );
  NAND2_X0P5A_A12TL \U1/U417  ( .A(\U1/rkey [26]), .B(\U1/n7 ), .Y(\U1/n309 )
         );
  AOI22_X0P5M_A12TL \U1/U416  ( .A0(\U1/key [26]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [26]), .B1(\U1/n1101 ), .Y(\U1/n310 ) );
  OAI211_X0P5M_A12TL \U1/U415  ( .A0(\U1/n1106 ), .A1(\U1/n308 ), .B0(
        \U1/n309 ), .C0(\U1/n310 ), .Y(\U1/n775 ) );
  INV_X0P5B_A12TL \U1/U414  ( .A(Kin[27]), .Y(\U1/n305 ) );
  NAND2_X0P5A_A12TL \U1/U413  ( .A(\U1/rkey [27]), .B(\U1/n7 ), .Y(\U1/n306 )
         );
  AOI22_X0P5M_A12TL \U1/U412  ( .A0(\U1/key [27]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [27]), .B1(\U1/n1101 ), .Y(\U1/n307 ) );
  OAI211_X0P5M_A12TL \U1/U411  ( .A0(\U1/n1106 ), .A1(\U1/n305 ), .B0(
        \U1/n306 ), .C0(\U1/n307 ), .Y(\U1/n774 ) );
  INV_X0P5B_A12TL \U1/U410  ( .A(Kin[28]), .Y(\U1/n302 ) );
  NAND2_X0P5A_A12TL \U1/U409  ( .A(\U1/rkey [28]), .B(\U1/n7 ), .Y(\U1/n303 )
         );
  AOI22_X0P5M_A12TL \U1/U408  ( .A0(\U1/key [28]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [28]), .B1(\U1/n1101 ), .Y(\U1/n304 ) );
  OAI211_X0P5M_A12TL \U1/U407  ( .A0(\U1/n1106 ), .A1(\U1/n302 ), .B0(
        \U1/n303 ), .C0(\U1/n304 ), .Y(\U1/n773 ) );
  INV_X0P5B_A12TL \U1/U406  ( .A(Kin[29]), .Y(\U1/n299 ) );
  NAND2_X0P5A_A12TL \U1/U405  ( .A(\U1/rkey [29]), .B(\U1/n7 ), .Y(\U1/n300 )
         );
  AOI22_X0P5M_A12TL \U1/U404  ( .A0(\U1/key [29]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [29]), .B1(\U1/n1101 ), .Y(\U1/n301 ) );
  OAI211_X0P5M_A12TL \U1/U403  ( .A0(\U1/n1106 ), .A1(\U1/n299 ), .B0(
        \U1/n300 ), .C0(\U1/n301 ), .Y(\U1/n772 ) );
  INV_X0P5B_A12TL \U1/U402  ( .A(Kin[30]), .Y(\U1/n296 ) );
  NAND2_X0P5A_A12TL \U1/U401  ( .A(\U1/rkey [30]), .B(\U1/n7 ), .Y(\U1/n297 )
         );
  AOI22_X0P5M_A12TL \U1/U400  ( .A0(\U1/key [30]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [30]), .B1(\U1/n1101 ), .Y(\U1/n298 ) );
  OAI211_X0P5M_A12TL \U1/U399  ( .A0(\U1/n1106 ), .A1(\U1/n296 ), .B0(
        \U1/n297 ), .C0(\U1/n298 ), .Y(\U1/n771 ) );
  INV_X0P5B_A12TL \U1/U398  ( .A(Kin[31]), .Y(\U1/n293 ) );
  NAND2_X0P5A_A12TL \U1/U397  ( .A(\U1/rkey [31]), .B(\U1/n7 ), .Y(\U1/n294 )
         );
  AOI22_X0P5M_A12TL \U1/U396  ( .A0(\U1/key [31]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [31]), .B1(\U1/n1101 ), .Y(\U1/n295 ) );
  OAI211_X0P5M_A12TL \U1/U395  ( .A0(\U1/n1106 ), .A1(\U1/n293 ), .B0(
        \U1/n294 ), .C0(\U1/n295 ), .Y(\U1/n770 ) );
  INV_X0P5B_A12TL \U1/U394  ( .A(Kin[32]), .Y(\U1/n290 ) );
  NAND2_X0P5A_A12TL \U1/U393  ( .A(\U1/rkey [32]), .B(\U1/n1099 ), .Y(
        \U1/n291 ) );
  AOI22_X0P5M_A12TL \U1/U392  ( .A0(\U1/key [32]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [32]), .B1(\U1/n1101 ), .Y(\U1/n292 ) );
  OAI211_X0P5M_A12TL \U1/U391  ( .A0(\U1/n1107 ), .A1(\U1/n290 ), .B0(
        \U1/n291 ), .C0(\U1/n292 ), .Y(\U1/n769 ) );
  INV_X0P5B_A12TL \U1/U390  ( .A(Kin[33]), .Y(\U1/n287 ) );
  NAND2_X0P5A_A12TL \U1/U389  ( .A(\U1/rkey [33]), .B(\U1/n7 ), .Y(\U1/n288 )
         );
  AOI22_X0P5M_A12TL \U1/U388  ( .A0(\U1/key [33]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [33]), .B1(\U1/n1101 ), .Y(\U1/n289 ) );
  OAI211_X0P5M_A12TL \U1/U387  ( .A0(\U1/n1105 ), .A1(\U1/n287 ), .B0(
        \U1/n288 ), .C0(\U1/n289 ), .Y(\U1/n768 ) );
  INV_X0P5B_A12TL \U1/U386  ( .A(Kin[34]), .Y(\U1/n284 ) );
  NAND2_X0P5A_A12TL \U1/U385  ( .A(\U1/rkey [34]), .B(\U1/n7 ), .Y(\U1/n285 )
         );
  AOI22_X0P5M_A12TL \U1/U384  ( .A0(\U1/key [34]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [34]), .B1(\U1/n1101 ), .Y(\U1/n286 ) );
  OAI211_X0P5M_A12TL \U1/U383  ( .A0(\U1/n1106 ), .A1(\U1/n284 ), .B0(
        \U1/n285 ), .C0(\U1/n286 ), .Y(\U1/n767 ) );
  INV_X0P5B_A12TL \U1/U382  ( .A(Kin[35]), .Y(\U1/n281 ) );
  NAND2_X0P5A_A12TL \U1/U381  ( .A(\U1/rkey [35]), .B(\U1/n7 ), .Y(\U1/n282 )
         );
  AOI22_X0P5M_A12TL \U1/U380  ( .A0(\U1/key [35]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [35]), .B1(\U1/n1100 ), .Y(\U1/n283 ) );
  OAI211_X0P5M_A12TL \U1/U379  ( .A0(\U1/n1104 ), .A1(\U1/n281 ), .B0(
        \U1/n282 ), .C0(\U1/n283 ), .Y(\U1/n766 ) );
  INV_X0P5B_A12TL \U1/U378  ( .A(Kin[36]), .Y(\U1/n278 ) );
  NAND2_X0P5A_A12TL \U1/U377  ( .A(\U1/rkey [36]), .B(\U1/n1099 ), .Y(
        \U1/n279 ) );
  AOI22_X0P5M_A12TL \U1/U376  ( .A0(\U1/key [36]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [36]), .B1(\U1/n1101 ), .Y(\U1/n280 ) );
  OAI211_X0P5M_A12TL \U1/U375  ( .A0(\U1/n1107 ), .A1(\U1/n278 ), .B0(
        \U1/n279 ), .C0(\U1/n280 ), .Y(\U1/n765 ) );
  INV_X0P5B_A12TL \U1/U374  ( .A(Kin[37]), .Y(\U1/n275 ) );
  NAND2_X0P5A_A12TL \U1/U373  ( .A(\U1/rkey [37]), .B(\U1/n1099 ), .Y(
        \U1/n276 ) );
  AOI22_X0P5M_A12TL \U1/U372  ( .A0(\U1/key [37]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [37]), .B1(\U1/n1100 ), .Y(\U1/n277 ) );
  OAI211_X0P5M_A12TL \U1/U371  ( .A0(\U1/n1106 ), .A1(\U1/n275 ), .B0(
        \U1/n276 ), .C0(\U1/n277 ), .Y(\U1/n764 ) );
  INV_X0P5B_A12TL \U1/U370  ( .A(Kin[38]), .Y(\U1/n272 ) );
  NAND2_X0P5A_A12TL \U1/U369  ( .A(\U1/rkey [38]), .B(\U1/n1099 ), .Y(
        \U1/n273 ) );
  AOI22_X0P5M_A12TL \U1/U368  ( .A0(\U1/key [38]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [38]), .B1(\U1/n1101 ), .Y(\U1/n274 ) );
  OAI211_X0P5M_A12TL \U1/U367  ( .A0(\U1/n1107 ), .A1(\U1/n272 ), .B0(
        \U1/n273 ), .C0(\U1/n274 ), .Y(\U1/n763 ) );
  INV_X0P5B_A12TL \U1/U366  ( .A(Kin[39]), .Y(\U1/n269 ) );
  NAND2_X0P5A_A12TL \U1/U365  ( .A(\U1/rkey [39]), .B(\U1/n1099 ), .Y(
        \U1/n270 ) );
  AOI22_X0P5M_A12TL \U1/U364  ( .A0(\U1/key [39]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [39]), .B1(\U1/n1101 ), .Y(\U1/n271 ) );
  OAI211_X0P5M_A12TL \U1/U363  ( .A0(\U1/n1105 ), .A1(\U1/n269 ), .B0(
        \U1/n270 ), .C0(\U1/n271 ), .Y(\U1/n762 ) );
  INV_X0P5B_A12TL \U1/U362  ( .A(Kin[40]), .Y(\U1/n266 ) );
  NAND2_X0P5A_A12TL \U1/U361  ( .A(\U1/rkey [40]), .B(\U1/n1099 ), .Y(
        \U1/n267 ) );
  AOI22_X0P5M_A12TL \U1/U360  ( .A0(\U1/key [40]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [40]), .B1(\U1/n1101 ), .Y(\U1/n268 ) );
  OAI211_X0P5M_A12TL \U1/U359  ( .A0(\U1/n1104 ), .A1(\U1/n266 ), .B0(
        \U1/n267 ), .C0(\U1/n268 ), .Y(\U1/n761 ) );
  INV_X0P5B_A12TL \U1/U358  ( .A(Kin[41]), .Y(\U1/n263 ) );
  NAND2_X0P5A_A12TL \U1/U357  ( .A(\U1/rkey [41]), .B(\U1/n1099 ), .Y(
        \U1/n264 ) );
  AOI22_X0P5M_A12TL \U1/U356  ( .A0(\U1/key [41]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [41]), .B1(\U1/n1101 ), .Y(\U1/n265 ) );
  OAI211_X0P5M_A12TL \U1/U355  ( .A0(\U1/n1106 ), .A1(\U1/n263 ), .B0(
        \U1/n264 ), .C0(\U1/n265 ), .Y(\U1/n760 ) );
  INV_X0P5B_A12TL \U1/U354  ( .A(Kin[42]), .Y(\U1/n260 ) );
  NAND2_X0P5A_A12TL \U1/U353  ( .A(\U1/rkey [42]), .B(\U1/n1099 ), .Y(
        \U1/n261 ) );
  AOI22_X0P5M_A12TL \U1/U352  ( .A0(\U1/key [42]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [42]), .B1(\U1/n1101 ), .Y(\U1/n262 ) );
  OAI211_X0P5M_A12TL \U1/U351  ( .A0(\U1/n1105 ), .A1(\U1/n260 ), .B0(
        \U1/n261 ), .C0(\U1/n262 ), .Y(\U1/n759 ) );
  INV_X0P5B_A12TL \U1/U350  ( .A(Kin[43]), .Y(\U1/n257 ) );
  NAND2_X0P5A_A12TL \U1/U349  ( .A(\U1/rkey [43]), .B(\U1/n1099 ), .Y(
        \U1/n258 ) );
  AOI22_X0P5M_A12TL \U1/U348  ( .A0(\U1/key [43]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [43]), .B1(\U1/n1101 ), .Y(\U1/n259 ) );
  OAI211_X0P5M_A12TL \U1/U347  ( .A0(\U1/n1104 ), .A1(\U1/n257 ), .B0(
        \U1/n258 ), .C0(\U1/n259 ), .Y(\U1/n758 ) );
  INV_X0P5B_A12TL \U1/U346  ( .A(Kin[44]), .Y(\U1/n254 ) );
  NAND2_X0P5A_A12TL \U1/U345  ( .A(\U1/rkey [44]), .B(\U1/n1099 ), .Y(
        \U1/n255 ) );
  AOI22_X0P5M_A12TL \U1/U344  ( .A0(\U1/key [44]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [44]), .B1(\U1/n1101 ), .Y(\U1/n256 ) );
  OAI211_X0P5M_A12TL \U1/U343  ( .A0(\U1/n1107 ), .A1(\U1/n254 ), .B0(
        \U1/n255 ), .C0(\U1/n256 ), .Y(\U1/n757 ) );
  INV_X0P5B_A12TL \U1/U342  ( .A(Kin[45]), .Y(\U1/n251 ) );
  NAND2_X0P5A_A12TL \U1/U341  ( .A(\U1/rkey [45]), .B(\U1/n1099 ), .Y(
        \U1/n252 ) );
  AOI22_X0P5M_A12TL \U1/U340  ( .A0(\U1/key [45]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [45]), .B1(\U1/n1101 ), .Y(\U1/n253 ) );
  OAI211_X0P5M_A12TL \U1/U339  ( .A0(\U1/n1105 ), .A1(\U1/n251 ), .B0(
        \U1/n252 ), .C0(\U1/n253 ), .Y(\U1/n756 ) );
  INV_X0P5B_A12TL \U1/U338  ( .A(Kin[46]), .Y(\U1/n248 ) );
  NAND2_X0P5A_A12TL \U1/U337  ( .A(\U1/rkey [46]), .B(\U1/n1099 ), .Y(
        \U1/n249 ) );
  AOI22_X0P5M_A12TL \U1/U336  ( .A0(\U1/key [46]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [46]), .B1(\U1/n1101 ), .Y(\U1/n250 ) );
  OAI211_X0P5M_A12TL \U1/U335  ( .A0(\U1/n1106 ), .A1(\U1/n248 ), .B0(
        \U1/n249 ), .C0(\U1/n250 ), .Y(\U1/n755 ) );
  INV_X0P5B_A12TL \U1/U334  ( .A(Kin[47]), .Y(\U1/n245 ) );
  NAND2_X0P5A_A12TL \U1/U333  ( .A(\U1/rkey [47]), .B(\U1/n1099 ), .Y(
        \U1/n246 ) );
  AOI22_X0P5M_A12TL \U1/U332  ( .A0(\U1/key [47]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [47]), .B1(\U1/n1101 ), .Y(\U1/n247 ) );
  OAI211_X0P5M_A12TL \U1/U331  ( .A0(\U1/n1106 ), .A1(\U1/n245 ), .B0(
        \U1/n246 ), .C0(\U1/n247 ), .Y(\U1/n754 ) );
  INV_X0P5B_A12TL \U1/U330  ( .A(Kin[48]), .Y(\U1/n242 ) );
  NAND2_X0P5A_A12TL \U1/U329  ( .A(\U1/rkey [48]), .B(\U1/n1099 ), .Y(
        \U1/n243 ) );
  AOI22_X0P5M_A12TL \U1/U328  ( .A0(\U1/key [48]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [48]), .B1(\U1/n1101 ), .Y(\U1/n244 ) );
  OAI211_X0P5M_A12TL \U1/U327  ( .A0(\U1/n1104 ), .A1(\U1/n242 ), .B0(
        \U1/n243 ), .C0(\U1/n244 ), .Y(\U1/n753 ) );
  INV_X0P5B_A12TL \U1/U326  ( .A(Kin[49]), .Y(\U1/n239 ) );
  NAND2_X0P5A_A12TL \U1/U325  ( .A(\U1/rkey [49]), .B(\U1/n1099 ), .Y(
        \U1/n240 ) );
  AOI22_X0P5M_A12TL \U1/U324  ( .A0(\U1/key [49]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [49]), .B1(\U1/n1101 ), .Y(\U1/n241 ) );
  OAI211_X0P5M_A12TL \U1/U323  ( .A0(\U1/n1104 ), .A1(\U1/n239 ), .B0(
        \U1/n240 ), .C0(\U1/n241 ), .Y(\U1/n752 ) );
  INV_X0P5B_A12TL \U1/U322  ( .A(Kin[50]), .Y(\U1/n236 ) );
  NAND2_X0P5A_A12TL \U1/U321  ( .A(\U1/rkey [50]), .B(\U1/n7 ), .Y(\U1/n237 )
         );
  AOI22_X0P5M_A12TL \U1/U320  ( .A0(\U1/key [50]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [50]), .B1(\U1/n1101 ), .Y(\U1/n238 ) );
  OAI211_X0P5M_A12TL \U1/U319  ( .A0(\U1/n1107 ), .A1(\U1/n236 ), .B0(
        \U1/n237 ), .C0(\U1/n238 ), .Y(\U1/n751 ) );
  INV_X0P5B_A12TL \U1/U318  ( .A(Kin[51]), .Y(\U1/n233 ) );
  NAND2_X0P5A_A12TL \U1/U317  ( .A(\U1/rkey [51]), .B(\U1/n1099 ), .Y(
        \U1/n234 ) );
  AOI22_X0P5M_A12TL \U1/U316  ( .A0(\U1/key [51]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [51]), .B1(\U1/n1101 ), .Y(\U1/n235 ) );
  OAI211_X0P5M_A12TL \U1/U315  ( .A0(\U1/n1104 ), .A1(\U1/n233 ), .B0(
        \U1/n234 ), .C0(\U1/n235 ), .Y(\U1/n750 ) );
  INV_X0P5B_A12TL \U1/U314  ( .A(Kin[52]), .Y(\U1/n230 ) );
  NAND2_X0P5A_A12TL \U1/U313  ( .A(\U1/rkey [52]), .B(\U1/n1099 ), .Y(
        \U1/n231 ) );
  AOI22_X0P5M_A12TL \U1/U312  ( .A0(\U1/key [52]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [52]), .B1(\U1/n1100 ), .Y(\U1/n232 ) );
  OAI211_X0P5M_A12TL \U1/U311  ( .A0(\U1/n1104 ), .A1(\U1/n230 ), .B0(
        \U1/n231 ), .C0(\U1/n232 ), .Y(\U1/n749 ) );
  INV_X0P5B_A12TL \U1/U310  ( .A(Kin[53]), .Y(\U1/n227 ) );
  NAND2_X0P5A_A12TL \U1/U309  ( .A(\U1/rkey [53]), .B(\U1/n1099 ), .Y(
        \U1/n228 ) );
  AOI22_X0P5M_A12TL \U1/U308  ( .A0(\U1/key [53]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [53]), .B1(\U1/n1100 ), .Y(\U1/n229 ) );
  OAI211_X0P5M_A12TL \U1/U307  ( .A0(\U1/n1104 ), .A1(\U1/n227 ), .B0(
        \U1/n228 ), .C0(\U1/n229 ), .Y(\U1/n748 ) );
  INV_X0P5B_A12TL \U1/U306  ( .A(Kin[54]), .Y(\U1/n224 ) );
  NAND2_X0P5A_A12TL \U1/U305  ( .A(\U1/rkey [54]), .B(\U1/n1099 ), .Y(
        \U1/n225 ) );
  AOI22_X0P5M_A12TL \U1/U304  ( .A0(\U1/key [54]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [54]), .B1(\U1/n1100 ), .Y(\U1/n226 ) );
  OAI211_X0P5M_A12TL \U1/U303  ( .A0(\U1/n1107 ), .A1(\U1/n224 ), .B0(
        \U1/n225 ), .C0(\U1/n226 ), .Y(\U1/n747 ) );
  INV_X0P5B_A12TL \U1/U302  ( .A(Kin[55]), .Y(\U1/n221 ) );
  NAND2_X0P5A_A12TL \U1/U301  ( .A(\U1/rkey [55]), .B(\U1/n1099 ), .Y(
        \U1/n222 ) );
  AOI22_X0P5M_A12TL \U1/U300  ( .A0(\U1/key [55]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [55]), .B1(\U1/n1100 ), .Y(\U1/n223 ) );
  OAI211_X0P5M_A12TL \U1/U299  ( .A0(\U1/n1105 ), .A1(\U1/n221 ), .B0(
        \U1/n222 ), .C0(\U1/n223 ), .Y(\U1/n746 ) );
  INV_X0P5B_A12TL \U1/U298  ( .A(Kin[56]), .Y(\U1/n218 ) );
  NAND2_X0P5A_A12TL \U1/U297  ( .A(\U1/rkey [56]), .B(\U1/n1099 ), .Y(
        \U1/n219 ) );
  AOI22_X0P5M_A12TL \U1/U296  ( .A0(\U1/key [56]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [56]), .B1(\U1/n1100 ), .Y(\U1/n220 ) );
  OAI211_X0P5M_A12TL \U1/U295  ( .A0(\U1/n1107 ), .A1(\U1/n218 ), .B0(
        \U1/n219 ), .C0(\U1/n220 ), .Y(\U1/n745 ) );
  INV_X0P5B_A12TL \U1/U294  ( .A(Kin[57]), .Y(\U1/n215 ) );
  NAND2_X0P5A_A12TL \U1/U293  ( .A(\U1/rkey [57]), .B(\U1/n1099 ), .Y(
        \U1/n216 ) );
  AOI22_X0P5M_A12TL \U1/U292  ( .A0(\U1/key [57]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [57]), .B1(\U1/n1100 ), .Y(\U1/n217 ) );
  OAI211_X0P5M_A12TL \U1/U291  ( .A0(\U1/n1107 ), .A1(\U1/n215 ), .B0(
        \U1/n216 ), .C0(\U1/n217 ), .Y(\U1/n744 ) );
  INV_X0P5B_A12TL \U1/U290  ( .A(Kin[58]), .Y(\U1/n212 ) );
  NAND2_X0P5A_A12TL \U1/U289  ( .A(\U1/rkey [58]), .B(\U1/n1099 ), .Y(
        \U1/n213 ) );
  AOI22_X0P5M_A12TL \U1/U288  ( .A0(\U1/key [58]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [58]), .B1(\U1/n1100 ), .Y(\U1/n214 ) );
  OAI211_X0P5M_A12TL \U1/U287  ( .A0(\U1/n1106 ), .A1(\U1/n212 ), .B0(
        \U1/n213 ), .C0(\U1/n214 ), .Y(\U1/n743 ) );
  INV_X0P5B_A12TL \U1/U286  ( .A(Kin[59]), .Y(\U1/n209 ) );
  NAND2_X0P5A_A12TL \U1/U285  ( .A(\U1/rkey [59]), .B(\U1/n1099 ), .Y(
        \U1/n210 ) );
  AOI22_X0P5M_A12TL \U1/U284  ( .A0(\U1/key [59]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [59]), .B1(\U1/n1100 ), .Y(\U1/n211 ) );
  OAI211_X0P5M_A12TL \U1/U283  ( .A0(\U1/n1105 ), .A1(\U1/n209 ), .B0(
        \U1/n210 ), .C0(\U1/n211 ), .Y(\U1/n742 ) );
  INV_X0P5B_A12TL \U1/U282  ( .A(Kin[60]), .Y(\U1/n206 ) );
  NAND2_X0P5A_A12TL \U1/U281  ( .A(\U1/rkey [60]), .B(\U1/n1099 ), .Y(
        \U1/n207 ) );
  AOI22_X0P5M_A12TL \U1/U280  ( .A0(\U1/key [60]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [60]), .B1(\U1/n1100 ), .Y(\U1/n208 ) );
  OAI211_X0P5M_A12TL \U1/U279  ( .A0(\U1/n1105 ), .A1(\U1/n206 ), .B0(
        \U1/n207 ), .C0(\U1/n208 ), .Y(\U1/n741 ) );
  INV_X0P5B_A12TL \U1/U278  ( .A(Kin[61]), .Y(\U1/n203 ) );
  NAND2_X0P5A_A12TL \U1/U277  ( .A(\U1/rkey [61]), .B(\U1/n1099 ), .Y(
        \U1/n204 ) );
  AOI22_X0P5M_A12TL \U1/U276  ( .A0(\U1/key [61]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [61]), .B1(\U1/n1100 ), .Y(\U1/n205 ) );
  OAI211_X0P5M_A12TL \U1/U275  ( .A0(\U1/n1104 ), .A1(\U1/n203 ), .B0(
        \U1/n204 ), .C0(\U1/n205 ), .Y(\U1/n740 ) );
  INV_X0P5B_A12TL \U1/U274  ( .A(Kin[62]), .Y(\U1/n200 ) );
  NAND2_X0P5A_A12TL \U1/U273  ( .A(\U1/rkey [62]), .B(\U1/n1099 ), .Y(
        \U1/n201 ) );
  AOI22_X0P5M_A12TL \U1/U272  ( .A0(\U1/key [62]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [62]), .B1(\U1/n1100 ), .Y(\U1/n202 ) );
  OAI211_X0P5M_A12TL \U1/U271  ( .A0(\U1/n1105 ), .A1(\U1/n200 ), .B0(
        \U1/n201 ), .C0(\U1/n202 ), .Y(\U1/n739 ) );
  INV_X0P5B_A12TL \U1/U270  ( .A(Kin[63]), .Y(\U1/n197 ) );
  NAND2_X0P5A_A12TL \U1/U269  ( .A(\U1/rkey [63]), .B(\U1/n1099 ), .Y(
        \U1/n198 ) );
  AOI22_X0P5M_A12TL \U1/U268  ( .A0(\U1/key [63]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [63]), .B1(\U1/n1100 ), .Y(\U1/n199 ) );
  OAI211_X0P5M_A12TL \U1/U267  ( .A0(\U1/n1104 ), .A1(\U1/n197 ), .B0(
        \U1/n198 ), .C0(\U1/n199 ), .Y(\U1/n738 ) );
  INV_X0P5B_A12TL \U1/U266  ( .A(Kin[64]), .Y(\U1/n194 ) );
  NAND2_X0P5A_A12TL \U1/U265  ( .A(\U1/rkey [64]), .B(\U1/n1099 ), .Y(
        \U1/n195 ) );
  AOI22_X0P5M_A12TL \U1/U264  ( .A0(\U1/key [64]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [64]), .B1(\U1/n1100 ), .Y(\U1/n196 ) );
  OAI211_X0P5M_A12TL \U1/U263  ( .A0(\U1/n1106 ), .A1(\U1/n194 ), .B0(
        \U1/n195 ), .C0(\U1/n196 ), .Y(\U1/n737 ) );
  INV_X0P5B_A12TL \U1/U262  ( .A(Kin[65]), .Y(\U1/n191 ) );
  NAND2_X0P5A_A12TL \U1/U261  ( .A(\U1/rkey [65]), .B(\U1/n1099 ), .Y(
        \U1/n192 ) );
  AOI22_X0P5M_A12TL \U1/U260  ( .A0(\U1/key [65]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [65]), .B1(\U1/n6 ), .Y(\U1/n193 ) );
  OAI211_X0P5M_A12TL \U1/U259  ( .A0(\U1/n1107 ), .A1(\U1/n191 ), .B0(
        \U1/n192 ), .C0(\U1/n193 ), .Y(\U1/n736 ) );
  INV_X0P5B_A12TL \U1/U258  ( .A(Kin[66]), .Y(\U1/n188 ) );
  NAND2_X0P5A_A12TL \U1/U257  ( .A(\U1/rkey [66]), .B(\U1/n1099 ), .Y(
        \U1/n189 ) );
  AOI22_X0P5M_A12TL \U1/U256  ( .A0(\U1/key [66]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [66]), .B1(\U1/n1100 ), .Y(\U1/n190 ) );
  OAI211_X0P5M_A12TL \U1/U255  ( .A0(\U1/n1107 ), .A1(\U1/n188 ), .B0(
        \U1/n189 ), .C0(\U1/n190 ), .Y(\U1/n735 ) );
  INV_X0P5B_A12TL \U1/U254  ( .A(Kin[67]), .Y(\U1/n185 ) );
  NAND2_X0P5A_A12TL \U1/U253  ( .A(\U1/rkey [67]), .B(\U1/n1099 ), .Y(
        \U1/n186 ) );
  AOI22_X0P5M_A12TL \U1/U252  ( .A0(\U1/key [67]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [67]), .B1(\U1/n1101 ), .Y(\U1/n187 ) );
  OAI211_X0P5M_A12TL \U1/U251  ( .A0(\U1/n1105 ), .A1(\U1/n185 ), .B0(
        \U1/n186 ), .C0(\U1/n187 ), .Y(\U1/n734 ) );
  INV_X0P5B_A12TL \U1/U250  ( .A(Kin[68]), .Y(\U1/n182 ) );
  NAND2_X0P5A_A12TL \U1/U249  ( .A(\U1/rkey [68]), .B(\U1/n1099 ), .Y(
        \U1/n183 ) );
  AOI22_X0P5M_A12TL \U1/U248  ( .A0(\U1/key [68]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [68]), .B1(\U1/n1101 ), .Y(\U1/n184 ) );
  OAI211_X0P5M_A12TL \U1/U247  ( .A0(\U1/n1106 ), .A1(\U1/n182 ), .B0(
        \U1/n183 ), .C0(\U1/n184 ), .Y(\U1/n733 ) );
  INV_X0P5B_A12TL \U1/U246  ( .A(Kin[69]), .Y(\U1/n179 ) );
  NAND2_X0P5A_A12TL \U1/U245  ( .A(\U1/rkey [69]), .B(\U1/n1099 ), .Y(
        \U1/n180 ) );
  AOI22_X0P5M_A12TL \U1/U244  ( .A0(\U1/key [69]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [69]), .B1(\U1/n1101 ), .Y(\U1/n181 ) );
  OAI211_X0P5M_A12TL \U1/U243  ( .A0(\U1/n1106 ), .A1(\U1/n179 ), .B0(
        \U1/n180 ), .C0(\U1/n181 ), .Y(\U1/n732 ) );
  INV_X0P5B_A12TL \U1/U242  ( .A(Kin[70]), .Y(\U1/n176 ) );
  NAND2_X0P5A_A12TL \U1/U241  ( .A(\U1/rkey [70]), .B(\U1/n1099 ), .Y(
        \U1/n177 ) );
  AOI22_X0P5M_A12TL \U1/U240  ( .A0(\U1/key [70]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [70]), .B1(\U1/n6 ), .Y(\U1/n178 ) );
  OAI211_X0P5M_A12TL \U1/U239  ( .A0(\U1/n1107 ), .A1(\U1/n176 ), .B0(
        \U1/n177 ), .C0(\U1/n178 ), .Y(\U1/n731 ) );
  INV_X0P5B_A12TL \U1/U238  ( .A(Kin[71]), .Y(\U1/n173 ) );
  NAND2_X0P5A_A12TL \U1/U237  ( .A(\U1/rkey [71]), .B(\U1/n1099 ), .Y(
        \U1/n174 ) );
  AOI22_X0P5M_A12TL \U1/U236  ( .A0(\U1/key [71]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [71]), .B1(\U1/n1101 ), .Y(\U1/n175 ) );
  OAI211_X0P5M_A12TL \U1/U235  ( .A0(\U1/n1104 ), .A1(\U1/n173 ), .B0(
        \U1/n174 ), .C0(\U1/n175 ), .Y(\U1/n730 ) );
  INV_X0P5B_A12TL \U1/U234  ( .A(Kin[72]), .Y(\U1/n170 ) );
  NAND2_X0P5A_A12TL \U1/U233  ( .A(\U1/rkey [72]), .B(\U1/n1099 ), .Y(
        \U1/n171 ) );
  AOI22_X0P5M_A12TL \U1/U232  ( .A0(\U1/key [72]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [72]), .B1(\U1/n6 ), .Y(\U1/n172 ) );
  OAI211_X0P5M_A12TL \U1/U231  ( .A0(\U1/n1105 ), .A1(\U1/n170 ), .B0(
        \U1/n171 ), .C0(\U1/n172 ), .Y(\U1/n729 ) );
  INV_X0P5B_A12TL \U1/U230  ( .A(Kin[73]), .Y(\U1/n167 ) );
  NAND2_X0P5A_A12TL \U1/U229  ( .A(\U1/rkey [73]), .B(\U1/n1099 ), .Y(
        \U1/n168 ) );
  AOI22_X0P5M_A12TL \U1/U228  ( .A0(\U1/key [73]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [73]), .B1(\U1/n6 ), .Y(\U1/n169 ) );
  OAI211_X0P5M_A12TL \U1/U227  ( .A0(\U1/n1104 ), .A1(\U1/n167 ), .B0(
        \U1/n168 ), .C0(\U1/n169 ), .Y(\U1/n728 ) );
  INV_X0P5B_A12TL \U1/U226  ( .A(Kin[74]), .Y(\U1/n164 ) );
  NAND2_X0P5A_A12TL \U1/U225  ( .A(\U1/rkey [74]), .B(\U1/n1099 ), .Y(
        \U1/n165 ) );
  AOI22_X0P5M_A12TL \U1/U224  ( .A0(\U1/key [74]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [74]), .B1(\U1/n6 ), .Y(\U1/n166 ) );
  OAI211_X0P5M_A12TL \U1/U223  ( .A0(\U1/n1106 ), .A1(\U1/n164 ), .B0(
        \U1/n165 ), .C0(\U1/n166 ), .Y(\U1/n727 ) );
  INV_X0P5B_A12TL \U1/U222  ( .A(Kin[75]), .Y(\U1/n161 ) );
  NAND2_X0P5A_A12TL \U1/U221  ( .A(\U1/rkey [75]), .B(\U1/n1099 ), .Y(
        \U1/n162 ) );
  AOI22_X0P5M_A12TL \U1/U220  ( .A0(\U1/key [75]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [75]), .B1(\U1/n6 ), .Y(\U1/n163 ) );
  OAI211_X0P5M_A12TL \U1/U219  ( .A0(\U1/n1104 ), .A1(\U1/n161 ), .B0(
        \U1/n162 ), .C0(\U1/n163 ), .Y(\U1/n726 ) );
  INV_X0P5B_A12TL \U1/U218  ( .A(Kin[76]), .Y(\U1/n158 ) );
  NAND2_X0P5A_A12TL \U1/U217  ( .A(\U1/rkey [76]), .B(\U1/n1099 ), .Y(
        \U1/n159 ) );
  AOI22_X0P5M_A12TL \U1/U216  ( .A0(\U1/key [76]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [76]), .B1(\U1/n6 ), .Y(\U1/n160 ) );
  OAI211_X0P5M_A12TL \U1/U215  ( .A0(\U1/n1106 ), .A1(\U1/n158 ), .B0(
        \U1/n159 ), .C0(\U1/n160 ), .Y(\U1/n725 ) );
  INV_X0P5B_A12TL \U1/U214  ( .A(Kin[77]), .Y(\U1/n155 ) );
  NAND2_X0P5A_A12TL \U1/U213  ( .A(\U1/rkey [77]), .B(\U1/n1099 ), .Y(
        \U1/n156 ) );
  AOI22_X0P5M_A12TL \U1/U212  ( .A0(\U1/key [77]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [77]), .B1(\U1/n6 ), .Y(\U1/n157 ) );
  OAI211_X0P5M_A12TL \U1/U211  ( .A0(\U1/n1106 ), .A1(\U1/n155 ), .B0(
        \U1/n156 ), .C0(\U1/n157 ), .Y(\U1/n724 ) );
  INV_X0P5B_A12TL \U1/U210  ( .A(Kin[78]), .Y(\U1/n152 ) );
  NAND2_X0P5A_A12TL \U1/U209  ( .A(\U1/rkey [78]), .B(\U1/n1099 ), .Y(
        \U1/n153 ) );
  AOI22_X0P5M_A12TL \U1/U208  ( .A0(\U1/key [78]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [78]), .B1(\U1/n6 ), .Y(\U1/n154 ) );
  OAI211_X0P5M_A12TL \U1/U207  ( .A0(\U1/n1106 ), .A1(\U1/n152 ), .B0(
        \U1/n153 ), .C0(\U1/n154 ), .Y(\U1/n723 ) );
  INV_X0P5B_A12TL \U1/U206  ( .A(Kin[79]), .Y(\U1/n149 ) );
  NAND2_X0P5A_A12TL \U1/U205  ( .A(\U1/rkey [79]), .B(\U1/n1099 ), .Y(
        \U1/n150 ) );
  AOI22_X0P5M_A12TL \U1/U204  ( .A0(\U1/key [79]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [79]), .B1(\U1/n1101 ), .Y(\U1/n151 ) );
  OAI211_X0P5M_A12TL \U1/U203  ( .A0(\U1/n1105 ), .A1(\U1/n149 ), .B0(
        \U1/n150 ), .C0(\U1/n151 ), .Y(\U1/n722 ) );
  INV_X0P5B_A12TL \U1/U202  ( .A(Kin[80]), .Y(\U1/n146 ) );
  NAND2_X0P5A_A12TL \U1/U201  ( .A(\U1/rkey [80]), .B(\U1/n1099 ), .Y(
        \U1/n147 ) );
  AOI22_X0P5M_A12TL \U1/U200  ( .A0(\U1/key [80]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [80]), .B1(\U1/n6 ), .Y(\U1/n148 ) );
  OAI211_X0P5M_A12TL \U1/U199  ( .A0(\U1/n1107 ), .A1(\U1/n146 ), .B0(
        \U1/n147 ), .C0(\U1/n148 ), .Y(\U1/n721 ) );
  INV_X0P5B_A12TL \U1/U198  ( .A(Kin[81]), .Y(\U1/n143 ) );
  NAND2_X0P5A_A12TL \U1/U197  ( .A(\U1/rkey [81]), .B(\U1/n1099 ), .Y(
        \U1/n144 ) );
  AOI22_X0P5M_A12TL \U1/U196  ( .A0(\U1/key [81]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [81]), .B1(\U1/n1101 ), .Y(\U1/n145 ) );
  OAI211_X0P5M_A12TL \U1/U195  ( .A0(\U1/n1106 ), .A1(\U1/n143 ), .B0(
        \U1/n144 ), .C0(\U1/n145 ), .Y(\U1/n720 ) );
  INV_X0P5B_A12TL \U1/U194  ( .A(Kin[82]), .Y(\U1/n140 ) );
  NAND2_X0P5A_A12TL \U1/U193  ( .A(\U1/rkey [82]), .B(\U1/n1099 ), .Y(
        \U1/n141 ) );
  AOI22_X0P5M_A12TL \U1/U192  ( .A0(\U1/key [82]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [82]), .B1(\U1/n6 ), .Y(\U1/n142 ) );
  OAI211_X0P5M_A12TL \U1/U191  ( .A0(\U1/n1107 ), .A1(\U1/n140 ), .B0(
        \U1/n141 ), .C0(\U1/n142 ), .Y(\U1/n719 ) );
  INV_X0P5B_A12TL \U1/U190  ( .A(Kin[83]), .Y(\U1/n137 ) );
  NAND2_X0P5A_A12TL \U1/U189  ( .A(\U1/rkey [83]), .B(\U1/n1099 ), .Y(
        \U1/n138 ) );
  AOI22_X0P5M_A12TL \U1/U188  ( .A0(\U1/key [83]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [83]), .B1(\U1/n1101 ), .Y(\U1/n139 ) );
  OAI211_X0P5M_A12TL \U1/U187  ( .A0(\U1/n1104 ), .A1(\U1/n137 ), .B0(
        \U1/n138 ), .C0(\U1/n139 ), .Y(\U1/n718 ) );
  INV_X0P5B_A12TL \U1/U186  ( .A(Kin[84]), .Y(\U1/n134 ) );
  NAND2_X0P5A_A12TL \U1/U185  ( .A(\U1/rkey [84]), .B(\U1/n1099 ), .Y(
        \U1/n135 ) );
  AOI22_X0P5M_A12TL \U1/U184  ( .A0(\U1/key [84]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [84]), .B1(\U1/n1101 ), .Y(\U1/n136 ) );
  OAI211_X0P5M_A12TL \U1/U183  ( .A0(\U1/n1105 ), .A1(\U1/n134 ), .B0(
        \U1/n135 ), .C0(\U1/n136 ), .Y(\U1/n717 ) );
  INV_X0P5B_A12TL \U1/U182  ( .A(Kin[85]), .Y(\U1/n131 ) );
  NAND2_X0P5A_A12TL \U1/U181  ( .A(\U1/rkey [85]), .B(\U1/n1099 ), .Y(
        \U1/n132 ) );
  AOI22_X0P5M_A12TL \U1/U180  ( .A0(\U1/key [85]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [85]), .B1(\U1/n1101 ), .Y(\U1/n133 ) );
  OAI211_X0P5M_A12TL \U1/U179  ( .A0(\U1/n1105 ), .A1(\U1/n131 ), .B0(
        \U1/n132 ), .C0(\U1/n133 ), .Y(\U1/n716 ) );
  INV_X0P5B_A12TL \U1/U178  ( .A(Kin[86]), .Y(\U1/n128 ) );
  NAND2_X0P5A_A12TL \U1/U177  ( .A(\U1/rkey [86]), .B(\U1/n1099 ), .Y(
        \U1/n129 ) );
  AOI22_X0P5M_A12TL \U1/U176  ( .A0(\U1/key [86]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [86]), .B1(\U1/n1101 ), .Y(\U1/n130 ) );
  OAI211_X0P5M_A12TL \U1/U175  ( .A0(\U1/n1105 ), .A1(\U1/n128 ), .B0(
        \U1/n129 ), .C0(\U1/n130 ), .Y(\U1/n715 ) );
  INV_X0P5B_A12TL \U1/U174  ( .A(Kin[87]), .Y(\U1/n125 ) );
  NAND2_X0P5A_A12TL \U1/U173  ( .A(\U1/rkey [87]), .B(\U1/n1099 ), .Y(
        \U1/n126 ) );
  AOI22_X0P5M_A12TL \U1/U172  ( .A0(\U1/key [87]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [87]), .B1(\U1/n1101 ), .Y(\U1/n127 ) );
  OAI211_X0P5M_A12TL \U1/U171  ( .A0(\U1/n1106 ), .A1(\U1/n125 ), .B0(
        \U1/n126 ), .C0(\U1/n127 ), .Y(\U1/n714 ) );
  INV_X0P5B_A12TL \U1/U170  ( .A(Kin[88]), .Y(\U1/n122 ) );
  NAND2_X0P5A_A12TL \U1/U169  ( .A(\U1/rkey [88]), .B(\U1/n1099 ), .Y(
        \U1/n123 ) );
  AOI22_X0P5M_A12TL \U1/U168  ( .A0(\U1/key [88]), .A1(\U1/n5 ), .B0(
        \U1/rkey_next [88]), .B1(\U1/n6 ), .Y(\U1/n124 ) );
  OAI211_X0P5M_A12TL \U1/U167  ( .A0(\U1/n1107 ), .A1(\U1/n122 ), .B0(
        \U1/n123 ), .C0(\U1/n124 ), .Y(\U1/n713 ) );
  INV_X0P5B_A12TL \U1/U166  ( .A(Kin[89]), .Y(\U1/n119 ) );
  NAND2_X0P5A_A12TL \U1/U165  ( .A(\U1/rkey [89]), .B(\U1/n1099 ), .Y(
        \U1/n120 ) );
  AOI22_X0P5M_A12TL \U1/U164  ( .A0(\U1/key [89]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [89]), .B1(\U1/n1101 ), .Y(\U1/n121 ) );
  OAI211_X0P5M_A12TL \U1/U163  ( .A0(\U1/n1106 ), .A1(\U1/n119 ), .B0(
        \U1/n120 ), .C0(\U1/n121 ), .Y(\U1/n712 ) );
  INV_X0P5B_A12TL \U1/U162  ( .A(Kin[90]), .Y(\U1/n116 ) );
  NAND2_X0P5A_A12TL \U1/U161  ( .A(\U1/rkey [90]), .B(\U1/n1099 ), .Y(
        \U1/n117 ) );
  AOI22_X0P5M_A12TL \U1/U160  ( .A0(\U1/key [90]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [90]), .B1(\U1/n6 ), .Y(\U1/n118 ) );
  OAI211_X0P5M_A12TL \U1/U159  ( .A0(\U1/n1107 ), .A1(\U1/n116 ), .B0(
        \U1/n117 ), .C0(\U1/n118 ), .Y(\U1/n711 ) );
  INV_X0P5B_A12TL \U1/U158  ( .A(Kin[91]), .Y(\U1/n113 ) );
  NAND2_X0P5A_A12TL \U1/U157  ( .A(\U1/rkey [91]), .B(\U1/n1099 ), .Y(
        \U1/n114 ) );
  AOI22_X0P5M_A12TL \U1/U156  ( .A0(\U1/key [91]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [91]), .B1(\U1/n1101 ), .Y(\U1/n115 ) );
  OAI211_X0P5M_A12TL \U1/U155  ( .A0(\U1/n1107 ), .A1(\U1/n113 ), .B0(
        \U1/n114 ), .C0(\U1/n115 ), .Y(\U1/n710 ) );
  INV_X0P5B_A12TL \U1/U154  ( .A(Kin[92]), .Y(\U1/n110 ) );
  NAND2_X0P5A_A12TL \U1/U153  ( .A(\U1/rkey [92]), .B(\U1/n1099 ), .Y(
        \U1/n111 ) );
  AOI22_X0P5M_A12TL \U1/U152  ( .A0(\U1/key [92]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [92]), .B1(\U1/n1101 ), .Y(\U1/n112 ) );
  OAI211_X0P5M_A12TL \U1/U151  ( .A0(\U1/n1104 ), .A1(\U1/n110 ), .B0(
        \U1/n111 ), .C0(\U1/n112 ), .Y(\U1/n709 ) );
  INV_X0P5B_A12TL \U1/U150  ( .A(Kin[93]), .Y(\U1/n107 ) );
  NAND2_X0P5A_A12TL \U1/U149  ( .A(\U1/rkey [93]), .B(\U1/n1099 ), .Y(
        \U1/n108 ) );
  AOI22_X0P5M_A12TL \U1/U148  ( .A0(\U1/key [93]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [93]), .B1(\U1/n1101 ), .Y(\U1/n109 ) );
  OAI211_X0P5M_A12TL \U1/U147  ( .A0(\U1/n1105 ), .A1(\U1/n107 ), .B0(
        \U1/n108 ), .C0(\U1/n109 ), .Y(\U1/n708 ) );
  INV_X0P5B_A12TL \U1/U146  ( .A(Kin[94]), .Y(\U1/n104 ) );
  NAND2_X0P5A_A12TL \U1/U145  ( .A(\U1/rkey [94]), .B(\U1/n1099 ), .Y(
        \U1/n105 ) );
  AOI22_X0P5M_A12TL \U1/U144  ( .A0(\U1/key [94]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [94]), .B1(\U1/n1101 ), .Y(\U1/n106 ) );
  OAI211_X0P5M_A12TL \U1/U143  ( .A0(\U1/n1107 ), .A1(\U1/n104 ), .B0(
        \U1/n105 ), .C0(\U1/n106 ), .Y(\U1/n707 ) );
  INV_X0P5B_A12TL \U1/U142  ( .A(Kin[95]), .Y(\U1/n101 ) );
  NAND2_X0P5A_A12TL \U1/U141  ( .A(\U1/rkey [95]), .B(\U1/n1099 ), .Y(
        \U1/n102 ) );
  AOI22_X0P5M_A12TL \U1/U140  ( .A0(\U1/key [95]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [95]), .B1(\U1/n1101 ), .Y(\U1/n103 ) );
  OAI211_X0P5M_A12TL \U1/U139  ( .A0(\U1/n1105 ), .A1(\U1/n101 ), .B0(
        \U1/n102 ), .C0(\U1/n103 ), .Y(\U1/n706 ) );
  INV_X0P5B_A12TL \U1/U138  ( .A(Kin[96]), .Y(\U1/n98 ) );
  NAND2_X0P5A_A12TL \U1/U137  ( .A(\U1/rkey [96]), .B(\U1/n1099 ), .Y(\U1/n99 ) );
  AOI22_X0P5M_A12TL \U1/U136  ( .A0(\U1/key [96]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [96]), .B1(\U1/n1101 ), .Y(\U1/n100 ) );
  OAI211_X0P5M_A12TL \U1/U135  ( .A0(\U1/n1106 ), .A1(\U1/n98 ), .B0(\U1/n99 ), 
        .C0(\U1/n100 ), .Y(\U1/n705 ) );
  INV_X0P5B_A12TL \U1/U134  ( .A(Kin[97]), .Y(\U1/n95 ) );
  NAND2_X0P5A_A12TL \U1/U133  ( .A(\U1/rkey [97]), .B(\U1/n1099 ), .Y(\U1/n96 ) );
  AOI22_X0P5M_A12TL \U1/U132  ( .A0(\U1/key [97]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [97]), .B1(\U1/n1101 ), .Y(\U1/n97 ) );
  OAI211_X0P5M_A12TL \U1/U131  ( .A0(\U1/n1107 ), .A1(\U1/n95 ), .B0(\U1/n96 ), 
        .C0(\U1/n97 ), .Y(\U1/n704 ) );
  INV_X0P5B_A12TL \U1/U130  ( .A(Kin[98]), .Y(\U1/n92 ) );
  NAND2_X0P5A_A12TL \U1/U129  ( .A(\U1/rkey [98]), .B(\U1/n1099 ), .Y(\U1/n93 ) );
  AOI22_X0P5M_A12TL \U1/U128  ( .A0(\U1/key [98]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [98]), .B1(\U1/n1100 ), .Y(\U1/n94 ) );
  OAI211_X0P5M_A12TL \U1/U127  ( .A0(\U1/n1107 ), .A1(\U1/n92 ), .B0(\U1/n93 ), 
        .C0(\U1/n94 ), .Y(\U1/n703 ) );
  INV_X0P5B_A12TL \U1/U126  ( .A(Kin[99]), .Y(\U1/n89 ) );
  NAND2_X0P5A_A12TL \U1/U125  ( .A(\U1/rkey [99]), .B(\U1/n1099 ), .Y(\U1/n90 ) );
  AOI22_X0P5M_A12TL \U1/U124  ( .A0(\U1/key [99]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [99]), .B1(\U1/n1101 ), .Y(\U1/n91 ) );
  OAI211_X0P5M_A12TL \U1/U123  ( .A0(\U1/n1106 ), .A1(\U1/n89 ), .B0(\U1/n90 ), 
        .C0(\U1/n91 ), .Y(\U1/n702 ) );
  INV_X0P5B_A12TL \U1/U122  ( .A(Kin[100]), .Y(\U1/n86 ) );
  NAND2_X0P5A_A12TL \U1/U121  ( .A(\U1/rkey [100]), .B(\U1/n1099 ), .Y(
        \U1/n87 ) );
  AOI22_X0P5M_A12TL \U1/U120  ( .A0(\U1/key [100]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [100]), .B1(\U1/n1100 ), .Y(\U1/n88 ) );
  OAI211_X0P5M_A12TL \U1/U119  ( .A0(\U1/n1104 ), .A1(\U1/n86 ), .B0(\U1/n87 ), 
        .C0(\U1/n88 ), .Y(\U1/n701 ) );
  INV_X0P5B_A12TL \U1/U118  ( .A(Kin[101]), .Y(\U1/n83 ) );
  NAND2_X0P5A_A12TL \U1/U117  ( .A(\U1/rkey [101]), .B(\U1/n1099 ), .Y(
        \U1/n84 ) );
  AOI22_X0P5M_A12TL \U1/U116  ( .A0(\U1/key [101]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [101]), .B1(\U1/n1101 ), .Y(\U1/n85 ) );
  OAI211_X0P5M_A12TL \U1/U115  ( .A0(\U1/n1104 ), .A1(\U1/n83 ), .B0(\U1/n84 ), 
        .C0(\U1/n85 ), .Y(\U1/n700 ) );
  INV_X0P5B_A12TL \U1/U114  ( .A(Kin[102]), .Y(\U1/n80 ) );
  NAND2_X0P5A_A12TL \U1/U113  ( .A(\U1/rkey [102]), .B(\U1/n1099 ), .Y(
        \U1/n81 ) );
  AOI22_X0P5M_A12TL \U1/U112  ( .A0(\U1/key [102]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [102]), .B1(\U1/n1100 ), .Y(\U1/n82 ) );
  OAI211_X0P5M_A12TL \U1/U111  ( .A0(\U1/n1105 ), .A1(\U1/n80 ), .B0(\U1/n81 ), 
        .C0(\U1/n82 ), .Y(\U1/n699 ) );
  INV_X0P5B_A12TL \U1/U110  ( .A(Kin[103]), .Y(\U1/n77 ) );
  NAND2_X0P5A_A12TL \U1/U109  ( .A(\U1/rkey [103]), .B(\U1/n7 ), .Y(\U1/n78 )
         );
  AOI22_X0P5M_A12TL \U1/U108  ( .A0(\U1/key [103]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [103]), .B1(\U1/n1100 ), .Y(\U1/n79 ) );
  OAI211_X0P5M_A12TL \U1/U107  ( .A0(\U1/n1105 ), .A1(\U1/n77 ), .B0(\U1/n78 ), 
        .C0(\U1/n79 ), .Y(\U1/n698 ) );
  INV_X0P5B_A12TL \U1/U106  ( .A(Kin[104]), .Y(\U1/n74 ) );
  NAND2_X0P5A_A12TL \U1/U105  ( .A(\U1/rkey [104]), .B(\U1/n7 ), .Y(\U1/n75 )
         );
  AOI22_X0P5M_A12TL \U1/U104  ( .A0(\U1/key [104]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [104]), .B1(\U1/n1101 ), .Y(\U1/n76 ) );
  OAI211_X0P5M_A12TL \U1/U103  ( .A0(\U1/n1107 ), .A1(\U1/n74 ), .B0(\U1/n75 ), 
        .C0(\U1/n76 ), .Y(\U1/n697 ) );
  INV_X0P5B_A12TL \U1/U102  ( .A(Kin[105]), .Y(\U1/n71 ) );
  NAND2_X0P5A_A12TL \U1/U101  ( .A(\U1/rkey [105]), .B(\U1/n1099 ), .Y(
        \U1/n72 ) );
  AOI22_X0P5M_A12TL \U1/U100  ( .A0(\U1/key [105]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [105]), .B1(\U1/n1101 ), .Y(\U1/n73 ) );
  OAI211_X0P5M_A12TL \U1/U99  ( .A0(\U1/n1104 ), .A1(\U1/n71 ), .B0(\U1/n72 ), 
        .C0(\U1/n73 ), .Y(\U1/n696 ) );
  INV_X0P5B_A12TL \U1/U98  ( .A(Kin[106]), .Y(\U1/n68 ) );
  NAND2_X0P5A_A12TL \U1/U97  ( .A(\U1/rkey [106]), .B(\U1/n7 ), .Y(\U1/n69 )
         );
  AOI22_X0P5M_A12TL \U1/U96  ( .A0(\U1/key [106]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [106]), .B1(\U1/n1101 ), .Y(\U1/n70 ) );
  OAI211_X0P5M_A12TL \U1/U95  ( .A0(\U1/n1104 ), .A1(\U1/n68 ), .B0(\U1/n69 ), 
        .C0(\U1/n70 ), .Y(\U1/n695 ) );
  INV_X0P5B_A12TL \U1/U94  ( .A(Kin[107]), .Y(\U1/n65 ) );
  NAND2_X0P5A_A12TL \U1/U93  ( .A(\U1/rkey [107]), .B(\U1/n1099 ), .Y(\U1/n66 ) );
  AOI22_X0P5M_A12TL \U1/U92  ( .A0(\U1/key [107]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [107]), .B1(\U1/n1101 ), .Y(\U1/n67 ) );
  OAI211_X0P5M_A12TL \U1/U91  ( .A0(\U1/n1107 ), .A1(\U1/n65 ), .B0(\U1/n66 ), 
        .C0(\U1/n67 ), .Y(\U1/n694 ) );
  INV_X0P5B_A12TL \U1/U90  ( .A(Kin[108]), .Y(\U1/n62 ) );
  NAND2_X0P5A_A12TL \U1/U89  ( .A(\U1/rkey [108]), .B(\U1/n7 ), .Y(\U1/n63 )
         );
  AOI22_X0P5M_A12TL \U1/U88  ( .A0(\U1/key [108]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [108]), .B1(\U1/n1100 ), .Y(\U1/n64 ) );
  OAI211_X0P5M_A12TL \U1/U87  ( .A0(\U1/n1106 ), .A1(\U1/n62 ), .B0(\U1/n63 ), 
        .C0(\U1/n64 ), .Y(\U1/n693 ) );
  INV_X0P5B_A12TL \U1/U86  ( .A(Kin[109]), .Y(\U1/n59 ) );
  NAND2_X0P5A_A12TL \U1/U85  ( .A(\U1/rkey [109]), .B(\U1/n1099 ), .Y(\U1/n60 ) );
  AOI22_X0P5M_A12TL \U1/U84  ( .A0(\U1/key [109]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [109]), .B1(\U1/n1100 ), .Y(\U1/n61 ) );
  OAI211_X0P5M_A12TL \U1/U83  ( .A0(\U1/n1105 ), .A1(\U1/n59 ), .B0(\U1/n60 ), 
        .C0(\U1/n61 ), .Y(\U1/n692 ) );
  INV_X0P5B_A12TL \U1/U82  ( .A(Kin[110]), .Y(\U1/n56 ) );
  NAND2_X0P5A_A12TL \U1/U81  ( .A(\U1/rkey [110]), .B(\U1/n7 ), .Y(\U1/n57 )
         );
  AOI22_X0P5M_A12TL \U1/U80  ( .A0(\U1/key [110]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [110]), .B1(\U1/n1100 ), .Y(\U1/n58 ) );
  OAI211_X0P5M_A12TL \U1/U79  ( .A0(\U1/n1106 ), .A1(\U1/n56 ), .B0(\U1/n57 ), 
        .C0(\U1/n58 ), .Y(\U1/n691 ) );
  INV_X0P5B_A12TL \U1/U78  ( .A(Kin[111]), .Y(\U1/n53 ) );
  NAND2_X0P5A_A12TL \U1/U77  ( .A(\U1/rkey [111]), .B(\U1/n1099 ), .Y(\U1/n54 ) );
  AOI22_X0P5M_A12TL \U1/U76  ( .A0(\U1/key [111]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [111]), .B1(\U1/n1100 ), .Y(\U1/n55 ) );
  OAI211_X0P5M_A12TL \U1/U75  ( .A0(\U1/n1105 ), .A1(\U1/n53 ), .B0(\U1/n54 ), 
        .C0(\U1/n55 ), .Y(\U1/n690 ) );
  INV_X0P5B_A12TL \U1/U74  ( .A(Kin[112]), .Y(\U1/n50 ) );
  NAND2_X0P5A_A12TL \U1/U73  ( .A(\U1/rkey [112]), .B(\U1/n7 ), .Y(\U1/n51 )
         );
  AOI22_X0P5M_A12TL \U1/U72  ( .A0(\U1/key [112]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [112]), .B1(\U1/n1100 ), .Y(\U1/n52 ) );
  OAI211_X0P5M_A12TL \U1/U71  ( .A0(\U1/n1106 ), .A1(\U1/n50 ), .B0(\U1/n51 ), 
        .C0(\U1/n52 ), .Y(\U1/n689 ) );
  INV_X0P5B_A12TL \U1/U70  ( .A(Kin[113]), .Y(\U1/n47 ) );
  NAND2_X0P5A_A12TL \U1/U69  ( .A(\U1/rkey [113]), .B(\U1/n1099 ), .Y(\U1/n48 ) );
  AOI22_X0P5M_A12TL \U1/U68  ( .A0(\U1/key [113]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [113]), .B1(\U1/n1100 ), .Y(\U1/n49 ) );
  OAI211_X0P5M_A12TL \U1/U67  ( .A0(\U1/n1107 ), .A1(\U1/n47 ), .B0(\U1/n48 ), 
        .C0(\U1/n49 ), .Y(\U1/n688 ) );
  INV_X0P5B_A12TL \U1/U66  ( .A(Kin[114]), .Y(\U1/n44 ) );
  NAND2_X0P5A_A12TL \U1/U65  ( .A(\U1/rkey [114]), .B(\U1/n7 ), .Y(\U1/n45 )
         );
  AOI22_X0P5M_A12TL \U1/U64  ( .A0(\U1/key [114]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [114]), .B1(\U1/n1100 ), .Y(\U1/n46 ) );
  OAI211_X0P5M_A12TL \U1/U63  ( .A0(\U1/n1104 ), .A1(\U1/n44 ), .B0(\U1/n45 ), 
        .C0(\U1/n46 ), .Y(\U1/n687 ) );
  INV_X0P5B_A12TL \U1/U62  ( .A(Kin[115]), .Y(\U1/n41 ) );
  NAND2_X0P5A_A12TL \U1/U61  ( .A(\U1/rkey [115]), .B(\U1/n7 ), .Y(\U1/n42 )
         );
  AOI22_X0P5M_A12TL \U1/U60  ( .A0(\U1/key [115]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [115]), .B1(\U1/n1100 ), .Y(\U1/n43 ) );
  OAI211_X0P5M_A12TL \U1/U59  ( .A0(\U1/n1106 ), .A1(\U1/n41 ), .B0(\U1/n42 ), 
        .C0(\U1/n43 ), .Y(\U1/n686 ) );
  INV_X0P5B_A12TL \U1/U58  ( .A(Kin[116]), .Y(\U1/n38 ) );
  NAND2_X0P5A_A12TL \U1/U57  ( .A(\U1/rkey [116]), .B(\U1/n7 ), .Y(\U1/n39 )
         );
  AOI22_X0P5M_A12TL \U1/U56  ( .A0(\U1/key [116]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [116]), .B1(\U1/n1100 ), .Y(\U1/n40 ) );
  OAI211_X0P5M_A12TL \U1/U55  ( .A0(\U1/n1105 ), .A1(\U1/n38 ), .B0(\U1/n39 ), 
        .C0(\U1/n40 ), .Y(\U1/n685 ) );
  INV_X0P5B_A12TL \U1/U54  ( .A(Kin[117]), .Y(\U1/n35 ) );
  NAND2_X0P5A_A12TL \U1/U53  ( .A(\U1/rkey [117]), .B(\U1/n1099 ), .Y(\U1/n36 ) );
  AOI22_X0P5M_A12TL \U1/U52  ( .A0(\U1/key [117]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [117]), .B1(\U1/n1101 ), .Y(\U1/n37 ) );
  OAI211_X0P5M_A12TL \U1/U51  ( .A0(\U1/n1107 ), .A1(\U1/n35 ), .B0(\U1/n36 ), 
        .C0(\U1/n37 ), .Y(\U1/n684 ) );
  INV_X0P5B_A12TL \U1/U50  ( .A(Kin[118]), .Y(\U1/n32 ) );
  NAND2_X0P5A_A12TL \U1/U49  ( .A(\U1/rkey [118]), .B(\U1/n7 ), .Y(\U1/n33 )
         );
  AOI22_X0P5M_A12TL \U1/U48  ( .A0(\U1/key [118]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [118]), .B1(\U1/n1100 ), .Y(\U1/n34 ) );
  OAI211_X0P5M_A12TL \U1/U47  ( .A0(\U1/n1106 ), .A1(\U1/n32 ), .B0(\U1/n33 ), 
        .C0(\U1/n34 ), .Y(\U1/n683 ) );
  INV_X0P5B_A12TL \U1/U46  ( .A(Kin[119]), .Y(\U1/n29 ) );
  NAND2_X0P5A_A12TL \U1/U45  ( .A(\U1/rkey [119]), .B(\U1/n7 ), .Y(\U1/n30 )
         );
  AOI22_X0P5M_A12TL \U1/U44  ( .A0(\U1/key [119]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [119]), .B1(\U1/n1100 ), .Y(\U1/n31 ) );
  OAI211_X0P5M_A12TL \U1/U43  ( .A0(\U1/n1104 ), .A1(\U1/n29 ), .B0(\U1/n30 ), 
        .C0(\U1/n31 ), .Y(\U1/n682 ) );
  INV_X0P5B_A12TL \U1/U42  ( .A(Kin[120]), .Y(\U1/n26 ) );
  NAND2_X0P5A_A12TL \U1/U41  ( .A(\U1/rkey [120]), .B(\U1/n7 ), .Y(\U1/n27 )
         );
  AOI22_X0P5M_A12TL \U1/U40  ( .A0(\U1/key [120]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [120]), .B1(\U1/n1101 ), .Y(\U1/n28 ) );
  OAI211_X0P5M_A12TL \U1/U39  ( .A0(\U1/n1106 ), .A1(\U1/n26 ), .B0(\U1/n27 ), 
        .C0(\U1/n28 ), .Y(\U1/n681 ) );
  INV_X0P5B_A12TL \U1/U38  ( .A(Kin[121]), .Y(\U1/n23 ) );
  NAND2_X0P5A_A12TL \U1/U37  ( .A(\U1/rkey [121]), .B(\U1/n7 ), .Y(\U1/n24 )
         );
  AOI22_X0P5M_A12TL \U1/U36  ( .A0(\U1/key [121]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [121]), .B1(\U1/n1101 ), .Y(\U1/n25 ) );
  OAI211_X0P5M_A12TL \U1/U35  ( .A0(\U1/n1107 ), .A1(\U1/n23 ), .B0(\U1/n24 ), 
        .C0(\U1/n25 ), .Y(\U1/n680 ) );
  INV_X0P5B_A12TL \U1/U34  ( .A(Kin[122]), .Y(\U1/n20 ) );
  NAND2_X0P5A_A12TL \U1/U33  ( .A(\U1/rkey [122]), .B(\U1/n7 ), .Y(\U1/n21 )
         );
  AOI22_X0P5M_A12TL \U1/U32  ( .A0(\U1/key [122]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [122]), .B1(\U1/n1101 ), .Y(\U1/n22 ) );
  OAI211_X0P5M_A12TL \U1/U31  ( .A0(\U1/n1107 ), .A1(\U1/n20 ), .B0(\U1/n21 ), 
        .C0(\U1/n22 ), .Y(\U1/n679 ) );
  INV_X0P5B_A12TL \U1/U30  ( .A(Kin[123]), .Y(\U1/n17 ) );
  NAND2_X0P5A_A12TL \U1/U29  ( .A(\U1/rkey [123]), .B(\U1/n7 ), .Y(\U1/n18 )
         );
  AOI22_X0P5M_A12TL \U1/U28  ( .A0(\U1/key [123]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [123]), .B1(\U1/n1101 ), .Y(\U1/n19 ) );
  OAI211_X0P5M_A12TL \U1/U27  ( .A0(\U1/n1107 ), .A1(\U1/n17 ), .B0(\U1/n18 ), 
        .C0(\U1/n19 ), .Y(\U1/n678 ) );
  INV_X0P5B_A12TL \U1/U26  ( .A(Kin[124]), .Y(\U1/n14 ) );
  NAND2_X0P5A_A12TL \U1/U25  ( .A(\U1/rkey [124]), .B(\U1/n1099 ), .Y(\U1/n15 ) );
  AOI22_X0P5M_A12TL \U1/U24  ( .A0(\U1/key [124]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [124]), .B1(\U1/n1101 ), .Y(\U1/n16 ) );
  OAI211_X0P5M_A12TL \U1/U23  ( .A0(\U1/n1104 ), .A1(\U1/n14 ), .B0(\U1/n15 ), 
        .C0(\U1/n16 ), .Y(\U1/n677 ) );
  INV_X0P5B_A12TL \U1/U22  ( .A(Kin[125]), .Y(\U1/n11 ) );
  NAND2_X0P5A_A12TL \U1/U21  ( .A(\U1/rkey [125]), .B(\U1/n1099 ), .Y(\U1/n12 ) );
  AOI22_X0P5M_A12TL \U1/U20  ( .A0(\U1/key [125]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [125]), .B1(\U1/n1101 ), .Y(\U1/n13 ) );
  OAI211_X0P5M_A12TL \U1/U19  ( .A0(\U1/n1107 ), .A1(\U1/n11 ), .B0(\U1/n12 ), 
        .C0(\U1/n13 ), .Y(\U1/n676 ) );
  INV_X0P5B_A12TL \U1/U18  ( .A(Kin[126]), .Y(\U1/n8 ) );
  NAND2_X0P5A_A12TL \U1/U17  ( .A(\U1/rkey [126]), .B(\U1/n7 ), .Y(\U1/n9 ) );
  AOI22_X0P5M_A12TL \U1/U16  ( .A0(\U1/key [126]), .A1(\U1/n1103 ), .B0(
        \U1/rkey_next [126]), .B1(\U1/n1101 ), .Y(\U1/n10 ) );
  OAI211_X0P5M_A12TL \U1/U15  ( .A0(\U1/n1107 ), .A1(\U1/n8 ), .B0(\U1/n9 ), 
        .C0(\U1/n10 ), .Y(\U1/n675 ) );
  INV_X0P5B_A12TL \U1/U14  ( .A(Kin[127]), .Y(\U1/n2 ) );
  NAND2_X0P5A_A12TL \U1/U13  ( .A(\U1/rkey [127]), .B(\U1/n1099 ), .Y(\U1/n3 )
         );
  AOI22_X0P5M_A12TL \U1/U12  ( .A0(\U1/key [127]), .A1(\U1/n1102 ), .B0(
        \U1/rkey_next [127]), .B1(\U1/n1101 ), .Y(\U1/n4 ) );
  OAI211_X0P5M_A12TL \U1/U11  ( .A0(\U1/n1105 ), .A1(\U1/n2 ), .B0(\U1/n3 ), 
        .C0(\U1/n4 ), .Y(\U1/n674 ) );
  INV_X0P5B_A12TL \U1/U10  ( .A(\U1/n808 ), .Y(\U1/rcon [0]) );
  INV_X0P5B_A12TL \U1/U9  ( .A(\U1/n807 ), .Y(\U1/rcon [1]) );
  INV_X0P5B_A12TL \U1/U8  ( .A(\U1/n806 ), .Y(\U1/rcon [2]) );
  INV_X0P5B_A12TL \U1/U7  ( .A(\U1/n805 ), .Y(\U1/rcon [3]) );
  INV_X0P5B_A12TL \U1/U6  ( .A(\U1/n804 ), .Y(\U1/rcon [4]) );
  INV_X0P5B_A12TL \U1/U5  ( .A(\U1/n803 ), .Y(\U1/rcon [5]) );
  INV_X0P5B_A12TL \U1/U4  ( .A(\U1/n802 ), .Y(\U1/rcon [6]) );
  BUFH_X1M_A12TL \U1/aes_core/U386  ( .A(\U1/aes_core/n2 ), .Y(
        \U1/aes_core/n258 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U385  ( .A(\U1/rkey_next [0]), .B(
        \U1/aes_core/sb2 [0]), .Y(\U1/aes_core/n256 ) );
  INV_X0P5B_A12TL \U1/aes_core/U384  ( .A(\U1/sel ), .Y(\U1/aes_core/n2 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U383  ( .A(\U1/rkey_next [0]), .B(
        \U1/aes_core/sc3 [0]), .Y(\U1/aes_core/n257 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U382  ( .A0(\U1/aes_core/n256 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n257 ), .Y(
        \U1/dat_next [0]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U381  ( .A(\U1/rkey_next [100]), .B(
        \U1/aes_core/sb3 [4]), .Y(\U1/aes_core/n254 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U380  ( .A(\U1/rkey_next [100]), .B(
        \U1/aes_core/sc0 [4]), .Y(\U1/aes_core/n255 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U379  ( .A0(\U1/aes_core/n254 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n255 ), .Y(
        \U1/dat_next [100]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U378  ( .A(\U1/rkey_next [101]), .B(
        \U1/aes_core/sb3 [5]), .Y(\U1/aes_core/n252 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U377  ( .A(\U1/rkey_next [101]), .B(
        \U1/aes_core/sc0 [5]), .Y(\U1/aes_core/n253 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U376  ( .A0(\U1/aes_core/n252 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n253 ), .Y(
        \U1/dat_next [101]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U375  ( .A(\U1/rkey_next [102]), .B(
        \U1/aes_core/sb3 [6]), .Y(\U1/aes_core/n250 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U374  ( .A(\U1/rkey_next [102]), .B(
        \U1/aes_core/sc0 [6]), .Y(\U1/aes_core/n251 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U373  ( .A0(\U1/aes_core/n250 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n251 ), .Y(
        \U1/dat_next [102]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U372  ( .A(\U1/rkey_next [103]), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/n248 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U371  ( .A(\U1/rkey_next [103]), .B(
        \U1/aes_core/sc0 [7]), .Y(\U1/aes_core/n249 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U370  ( .A0(\U1/aes_core/n248 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n249 ), .Y(
        \U1/dat_next [103]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U369  ( .A(\U1/rkey_next [104]), .B(
        \U1/aes_core/sb2 [8]), .Y(\U1/aes_core/n246 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U368  ( .A(\U1/rkey_next [104]), .B(
        \U1/aes_core/sc0 [8]), .Y(\U1/aes_core/n247 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U367  ( .A0(\U1/aes_core/n246 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n247 ), .Y(
        \U1/dat_next [104]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U366  ( .A(\U1/rkey_next [105]), .B(
        \U1/aes_core/sb2 [9]), .Y(\U1/aes_core/n244 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U365  ( .A(\U1/rkey_next [105]), .B(
        \U1/aes_core/sc0 [9]), .Y(\U1/aes_core/n245 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U364  ( .A0(\U1/aes_core/n244 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n245 ), .Y(
        \U1/dat_next [105]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U363  ( .A(\U1/rkey_next [106]), .B(
        \U1/aes_core/sb2 [10]), .Y(\U1/aes_core/n242 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U362  ( .A(\U1/rkey_next [106]), .B(
        \U1/aes_core/sc0 [10]), .Y(\U1/aes_core/n243 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U361  ( .A0(\U1/aes_core/n242 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n243 ), .Y(
        \U1/dat_next [106]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U360  ( .A(\U1/rkey_next [107]), .B(
        \U1/aes_core/sb2 [11]), .Y(\U1/aes_core/n240 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U359  ( .A(\U1/rkey_next [107]), .B(
        \U1/aes_core/sc0 [11]), .Y(\U1/aes_core/n241 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U358  ( .A0(\U1/aes_core/n240 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n241 ), .Y(
        \U1/dat_next [107]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U357  ( .A(\U1/rkey_next [108]), .B(
        \U1/aes_core/sb2 [12]), .Y(\U1/aes_core/n238 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U356  ( .A(\U1/rkey_next [108]), .B(
        \U1/aes_core/sc0 [12]), .Y(\U1/aes_core/n239 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U355  ( .A0(\U1/aes_core/n238 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n239 ), .Y(
        \U1/dat_next [108]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U354  ( .A(\U1/rkey_next [109]), .B(
        \U1/aes_core/sb2 [13]), .Y(\U1/aes_core/n236 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U353  ( .A(\U1/rkey_next [109]), .B(
        \U1/aes_core/sc0 [13]), .Y(\U1/aes_core/n237 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U352  ( .A0(\U1/aes_core/n236 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n237 ), .Y(
        \U1/dat_next [109]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U351  ( .A(\U1/rkey_next [10]), .B(
        \U1/aes_core/sb1 [10]), .Y(\U1/aes_core/n234 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U350  ( .A(\U1/rkey_next [10]), .B(
        \U1/aes_core/sc3 [10]), .Y(\U1/aes_core/n235 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U349  ( .A0(\U1/aes_core/n234 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n235 ), .Y(
        \U1/dat_next [10]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U348  ( .A(\U1/rkey_next [110]), .B(
        \U1/aes_core/sb2 [14]), .Y(\U1/aes_core/n232 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U347  ( .A(\U1/rkey_next [110]), .B(
        \U1/aes_core/sc0 [14]), .Y(\U1/aes_core/n233 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U346  ( .A0(\U1/aes_core/n232 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n233 ), .Y(
        \U1/dat_next [110]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U345  ( .A(\U1/rkey_next [111]), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/n230 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U344  ( .A(\U1/rkey_next [111]), .B(
        \U1/aes_core/sc0 [15]), .Y(\U1/aes_core/n231 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U343  ( .A0(\U1/aes_core/n230 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n231 ), .Y(
        \U1/dat_next [111]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U342  ( .A(\U1/rkey_next [112]), .B(
        \U1/aes_core/sb1 [16]), .Y(\U1/aes_core/n228 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U341  ( .A(\U1/rkey_next [112]), .B(
        \U1/aes_core/sc0 [16]), .Y(\U1/aes_core/n229 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U340  ( .A0(\U1/aes_core/n228 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n229 ), .Y(
        \U1/dat_next [112]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U339  ( .A(\U1/rkey_next [113]), .B(
        \U1/aes_core/sb1 [17]), .Y(\U1/aes_core/n226 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U338  ( .A(\U1/rkey_next [113]), .B(
        \U1/aes_core/sc0 [17]), .Y(\U1/aes_core/n227 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U337  ( .A0(\U1/aes_core/n226 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n227 ), .Y(
        \U1/dat_next [113]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U336  ( .A(\U1/rkey_next [114]), .B(
        \U1/aes_core/sb1 [18]), .Y(\U1/aes_core/n224 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U335  ( .A(\U1/rkey_next [114]), .B(
        \U1/aes_core/sc0 [18]), .Y(\U1/aes_core/n225 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U334  ( .A0(\U1/aes_core/n224 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n225 ), .Y(
        \U1/dat_next [114]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U333  ( .A(\U1/rkey_next [115]), .B(
        \U1/aes_core/sb1 [19]), .Y(\U1/aes_core/n222 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U332  ( .A(\U1/rkey_next [115]), .B(
        \U1/aes_core/sc0 [19]), .Y(\U1/aes_core/n223 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U331  ( .A0(\U1/aes_core/n222 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n223 ), .Y(
        \U1/dat_next [115]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U330  ( .A(\U1/rkey_next [116]), .B(
        \U1/aes_core/sb1 [20]), .Y(\U1/aes_core/n220 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U329  ( .A(\U1/rkey_next [116]), .B(
        \U1/aes_core/sc0 [20]), .Y(\U1/aes_core/n221 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U328  ( .A0(\U1/aes_core/n220 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n221 ), .Y(
        \U1/dat_next [116]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U327  ( .A(\U1/rkey_next [117]), .B(
        \U1/aes_core/sb1 [21]), .Y(\U1/aes_core/n218 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U326  ( .A(\U1/rkey_next [117]), .B(
        \U1/aes_core/sc0 [21]), .Y(\U1/aes_core/n219 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U325  ( .A0(\U1/aes_core/n218 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n219 ), .Y(
        \U1/dat_next [117]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U324  ( .A(\U1/rkey_next [118]), .B(
        \U1/aes_core/sb1 [22]), .Y(\U1/aes_core/n216 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U323  ( .A(\U1/rkey_next [118]), .B(
        \U1/aes_core/sc0 [22]), .Y(\U1/aes_core/n217 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U322  ( .A0(\U1/aes_core/n216 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n217 ), .Y(
        \U1/dat_next [118]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U321  ( .A(\U1/rkey_next [119]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/n214 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U320  ( .A(\U1/rkey_next [119]), .B(
        \U1/aes_core/sc0 [23]), .Y(\U1/aes_core/n215 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U319  ( .A0(\U1/aes_core/n214 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n215 ), .Y(
        \U1/dat_next [119]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U318  ( .A(\U1/rkey_next [11]), .B(
        \U1/aes_core/sb1 [11]), .Y(\U1/aes_core/n212 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U317  ( .A(\U1/rkey_next [11]), .B(
        \U1/aes_core/sc3 [11]), .Y(\U1/aes_core/n213 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U316  ( .A0(\U1/aes_core/n212 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n213 ), .Y(
        \U1/dat_next [11]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U315  ( .A(\U1/rkey_next [120]), .B(
        \U1/aes_core/sb0 [24]), .Y(\U1/aes_core/n210 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U314  ( .A(\U1/rkey_next [120]), .B(
        \U1/aes_core/sc0 [24]), .Y(\U1/aes_core/n211 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U313  ( .A0(\U1/aes_core/n210 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n211 ), .Y(
        \U1/dat_next [120]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U312  ( .A(\U1/rkey_next [121]), .B(
        \U1/aes_core/sb0 [25]), .Y(\U1/aes_core/n208 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U311  ( .A(\U1/rkey_next [121]), .B(
        \U1/aes_core/sc0 [25]), .Y(\U1/aes_core/n209 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U310  ( .A0(\U1/aes_core/n208 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n209 ), .Y(
        \U1/dat_next [121]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U309  ( .A(\U1/rkey_next [122]), .B(
        \U1/aes_core/sb0 [26]), .Y(\U1/aes_core/n206 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U308  ( .A(\U1/rkey_next [122]), .B(
        \U1/aes_core/sc0 [26]), .Y(\U1/aes_core/n207 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U307  ( .A0(\U1/aes_core/n206 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n207 ), .Y(
        \U1/dat_next [122]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U306  ( .A(\U1/rkey_next [123]), .B(
        \U1/aes_core/sb0 [27]), .Y(\U1/aes_core/n204 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U305  ( .A(\U1/rkey_next [123]), .B(
        \U1/aes_core/sc0 [27]), .Y(\U1/aes_core/n205 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U304  ( .A0(\U1/aes_core/n204 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n205 ), .Y(
        \U1/dat_next [123]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U303  ( .A(\U1/rkey_next [124]), .B(
        \U1/aes_core/sb0 [28]), .Y(\U1/aes_core/n202 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U302  ( .A(\U1/rkey_next [124]), .B(
        \U1/aes_core/sc0 [28]), .Y(\U1/aes_core/n203 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U301  ( .A0(\U1/aes_core/n202 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n203 ), .Y(
        \U1/dat_next [124]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U300  ( .A(\U1/rkey_next [125]), .B(
        \U1/aes_core/sb0 [29]), .Y(\U1/aes_core/n200 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U299  ( .A(\U1/rkey_next [125]), .B(
        \U1/aes_core/sc0 [29]), .Y(\U1/aes_core/n201 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U298  ( .A0(\U1/aes_core/n200 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n201 ), .Y(
        \U1/dat_next [125]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U297  ( .A(\U1/rkey_next [126]), .B(
        \U1/aes_core/sb0 [30]), .Y(\U1/aes_core/n198 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U296  ( .A(\U1/rkey_next [126]), .B(
        \U1/aes_core/sc0 [30]), .Y(\U1/aes_core/n199 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U295  ( .A0(\U1/aes_core/n198 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n199 ), .Y(
        \U1/dat_next [126]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U294  ( .A(\U1/rkey_next [127]), .B(
        \U1/aes_core/sb0 [31]), .Y(\U1/aes_core/n196 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U293  ( .A(\U1/rkey_next [127]), .B(
        \U1/aes_core/sc0 [31]), .Y(\U1/aes_core/n197 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U292  ( .A0(\U1/aes_core/n196 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n197 ), .Y(
        \U1/dat_next [127]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U291  ( .A(\U1/rkey_next [12]), .B(
        \U1/aes_core/sb1 [12]), .Y(\U1/aes_core/n194 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U290  ( .A(\U1/rkey_next [12]), .B(
        \U1/aes_core/sc3 [12]), .Y(\U1/aes_core/n195 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U289  ( .A0(\U1/aes_core/n194 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n195 ), .Y(
        \U1/dat_next [12]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U288  ( .A(\U1/rkey_next [13]), .B(
        \U1/aes_core/sb1 [13]), .Y(\U1/aes_core/n192 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U287  ( .A(\U1/rkey_next [13]), .B(
        \U1/aes_core/sc3 [13]), .Y(\U1/aes_core/n193 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U286  ( .A0(\U1/aes_core/n192 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n193 ), .Y(
        \U1/dat_next [13]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U285  ( .A(\U1/rkey_next [14]), .B(
        \U1/aes_core/sb1 [14]), .Y(\U1/aes_core/n190 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U284  ( .A(\U1/rkey_next [14]), .B(
        \U1/aes_core/sc3 [14]), .Y(\U1/aes_core/n191 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U283  ( .A0(\U1/aes_core/n190 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n191 ), .Y(
        \U1/dat_next [14]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U282  ( .A(\U1/rkey_next [15]), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/n188 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U281  ( .A(\U1/rkey_next [15]), .B(
        \U1/aes_core/sc3 [15]), .Y(\U1/aes_core/n189 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U280  ( .A0(\U1/aes_core/n188 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n189 ), .Y(
        \U1/dat_next [15]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U279  ( .A(\U1/rkey_next [16]), .B(
        \U1/aes_core/sb0 [16]), .Y(\U1/aes_core/n186 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U278  ( .A(\U1/rkey_next [16]), .B(
        \U1/aes_core/sc3 [16]), .Y(\U1/aes_core/n187 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U277  ( .A0(\U1/aes_core/n186 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n187 ), .Y(
        \U1/dat_next [16]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U276  ( .A(\U1/rkey_next [17]), .B(
        \U1/aes_core/sb0 [17]), .Y(\U1/aes_core/n184 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U275  ( .A(\U1/rkey_next [17]), .B(
        \U1/aes_core/sc3 [17]), .Y(\U1/aes_core/n185 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U274  ( .A0(\U1/aes_core/n184 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n185 ), .Y(
        \U1/dat_next [17]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U273  ( .A(\U1/rkey_next [18]), .B(
        \U1/aes_core/sb0 [18]), .Y(\U1/aes_core/n182 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U272  ( .A(\U1/rkey_next [18]), .B(
        \U1/aes_core/sc3 [18]), .Y(\U1/aes_core/n183 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U271  ( .A0(\U1/aes_core/n182 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n183 ), .Y(
        \U1/dat_next [18]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U270  ( .A(\U1/rkey_next [19]), .B(
        \U1/aes_core/sb0 [19]), .Y(\U1/aes_core/n180 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U269  ( .A(\U1/rkey_next [19]), .B(
        \U1/aes_core/sc3 [19]), .Y(\U1/aes_core/n181 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U268  ( .A0(\U1/aes_core/n180 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n181 ), .Y(
        \U1/dat_next [19]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U267  ( .A(\U1/rkey_next [1]), .B(
        \U1/aes_core/sb2 [1]), .Y(\U1/aes_core/n178 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U266  ( .A(\U1/rkey_next [1]), .B(
        \U1/aes_core/sc3 [1]), .Y(\U1/aes_core/n179 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U265  ( .A0(\U1/aes_core/n178 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n179 ), .Y(
        \U1/dat_next [1]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U264  ( .A(\U1/rkey_next [20]), .B(
        \U1/aes_core/sb0 [20]), .Y(\U1/aes_core/n176 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U263  ( .A(\U1/rkey_next [20]), .B(
        \U1/aes_core/sc3 [20]), .Y(\U1/aes_core/n177 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U262  ( .A0(\U1/aes_core/n176 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n177 ), .Y(
        \U1/dat_next [20]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U261  ( .A(\U1/rkey_next [21]), .B(
        \U1/aes_core/sb0 [21]), .Y(\U1/aes_core/n174 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U260  ( .A(\U1/rkey_next [21]), .B(
        \U1/aes_core/sc3 [21]), .Y(\U1/aes_core/n175 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U259  ( .A0(\U1/aes_core/n174 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n175 ), .Y(
        \U1/dat_next [21]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U258  ( .A(\U1/rkey_next [22]), .B(
        \U1/aes_core/sb0 [22]), .Y(\U1/aes_core/n172 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U257  ( .A(\U1/rkey_next [22]), .B(
        \U1/aes_core/sc3 [22]), .Y(\U1/aes_core/n173 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U256  ( .A0(\U1/aes_core/n172 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n173 ), .Y(
        \U1/dat_next [22]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U255  ( .A(\U1/rkey_next [23]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/n170 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U254  ( .A(\U1/rkey_next [23]), .B(
        \U1/aes_core/sc3 [23]), .Y(\U1/aes_core/n171 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U253  ( .A0(\U1/aes_core/n170 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n171 ), .Y(
        \U1/dat_next [23]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U252  ( .A(\U1/rkey_next [24]), .B(
        \U1/aes_core/sb3 [24]), .Y(\U1/aes_core/n168 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U251  ( .A(\U1/rkey_next [24]), .B(
        \U1/aes_core/sc3 [24]), .Y(\U1/aes_core/n169 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U250  ( .A0(\U1/aes_core/n168 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n169 ), .Y(
        \U1/dat_next [24]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U249  ( .A(\U1/rkey_next [25]), .B(
        \U1/aes_core/sb3 [25]), .Y(\U1/aes_core/n166 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U248  ( .A(\U1/rkey_next [25]), .B(
        \U1/aes_core/sc3 [25]), .Y(\U1/aes_core/n167 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U247  ( .A0(\U1/aes_core/n166 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n167 ), .Y(
        \U1/dat_next [25]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U246  ( .A(\U1/rkey_next [26]), .B(
        \U1/aes_core/sb3 [26]), .Y(\U1/aes_core/n164 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U245  ( .A(\U1/rkey_next [26]), .B(
        \U1/aes_core/sc3 [26]), .Y(\U1/aes_core/n165 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U244  ( .A0(\U1/aes_core/n164 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n165 ), .Y(
        \U1/dat_next [26]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U243  ( .A(\U1/rkey_next [27]), .B(
        \U1/aes_core/sb3 [27]), .Y(\U1/aes_core/n162 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U242  ( .A(\U1/rkey_next [27]), .B(
        \U1/aes_core/sc3 [27]), .Y(\U1/aes_core/n163 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U241  ( .A0(\U1/aes_core/n162 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n163 ), .Y(
        \U1/dat_next [27]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U240  ( .A(\U1/rkey_next [28]), .B(
        \U1/aes_core/sb3 [28]), .Y(\U1/aes_core/n160 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U239  ( .A(\U1/rkey_next [28]), .B(
        \U1/aes_core/sc3 [28]), .Y(\U1/aes_core/n161 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U238  ( .A0(\U1/aes_core/n160 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n161 ), .Y(
        \U1/dat_next [28]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U237  ( .A(\U1/rkey_next [29]), .B(
        \U1/aes_core/sb3 [29]), .Y(\U1/aes_core/n158 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U236  ( .A(\U1/rkey_next [29]), .B(
        \U1/aes_core/sc3 [29]), .Y(\U1/aes_core/n159 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U235  ( .A0(\U1/aes_core/n158 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n159 ), .Y(
        \U1/dat_next [29]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U234  ( .A(\U1/rkey_next [2]), .B(
        \U1/aes_core/sb2 [2]), .Y(\U1/aes_core/n156 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U233  ( .A(\U1/rkey_next [2]), .B(
        \U1/aes_core/sc3 [2]), .Y(\U1/aes_core/n157 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U232  ( .A0(\U1/aes_core/n156 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n157 ), .Y(
        \U1/dat_next [2]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U231  ( .A(\U1/rkey_next [30]), .B(
        \U1/aes_core/sb3 [30]), .Y(\U1/aes_core/n154 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U230  ( .A(\U1/rkey_next [30]), .B(
        \U1/aes_core/sc3 [30]), .Y(\U1/aes_core/n155 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U229  ( .A0(\U1/aes_core/n154 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n155 ), .Y(
        \U1/dat_next [30]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U228  ( .A(\U1/rkey_next [31]), .B(
        \U1/aes_core/sb3 [31]), .Y(\U1/aes_core/n152 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U227  ( .A(\U1/rkey_next [31]), .B(
        \U1/aes_core/sc3 [31]), .Y(\U1/aes_core/n153 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U226  ( .A0(\U1/aes_core/n152 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n153 ), .Y(
        \U1/dat_next [31]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U225  ( .A(\U1/rkey_next [32]), .B(
        \U1/aes_core/sb1 [0]), .Y(\U1/aes_core/n150 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U224  ( .A(\U1/rkey_next [32]), .B(
        \U1/aes_core/sc2 [0]), .Y(\U1/aes_core/n151 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U223  ( .A0(\U1/aes_core/n150 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n151 ), .Y(
        \U1/dat_next [32]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U222  ( .A(\U1/rkey_next [33]), .B(
        \U1/aes_core/sb1 [1]), .Y(\U1/aes_core/n148 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U221  ( .A(\U1/rkey_next [33]), .B(
        \U1/aes_core/sc2 [1]), .Y(\U1/aes_core/n149 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U220  ( .A0(\U1/aes_core/n148 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n149 ), .Y(
        \U1/dat_next [33]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U219  ( .A(\U1/rkey_next [34]), .B(
        \U1/aes_core/sb1 [2]), .Y(\U1/aes_core/n146 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U218  ( .A(\U1/rkey_next [34]), .B(
        \U1/aes_core/sc2 [2]), .Y(\U1/aes_core/n147 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U217  ( .A0(\U1/aes_core/n146 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n147 ), .Y(
        \U1/dat_next [34]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U216  ( .A(\U1/rkey_next [35]), .B(
        \U1/aes_core/sb1 [3]), .Y(\U1/aes_core/n144 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U215  ( .A(\U1/rkey_next [35]), .B(
        \U1/aes_core/sc2 [3]), .Y(\U1/aes_core/n145 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U214  ( .A0(\U1/aes_core/n144 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n145 ), .Y(
        \U1/dat_next [35]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U213  ( .A(\U1/rkey_next [36]), .B(
        \U1/aes_core/sb1 [4]), .Y(\U1/aes_core/n142 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U212  ( .A(\U1/rkey_next [36]), .B(
        \U1/aes_core/sc2 [4]), .Y(\U1/aes_core/n143 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U211  ( .A0(\U1/aes_core/n142 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n143 ), .Y(
        \U1/dat_next [36]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U210  ( .A(\U1/rkey_next [37]), .B(
        \U1/aes_core/sb1 [5]), .Y(\U1/aes_core/n140 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U209  ( .A(\U1/rkey_next [37]), .B(
        \U1/aes_core/sc2 [5]), .Y(\U1/aes_core/n141 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U208  ( .A0(\U1/aes_core/n140 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n141 ), .Y(
        \U1/dat_next [37]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U207  ( .A(\U1/rkey_next [38]), .B(
        \U1/aes_core/sb1 [6]), .Y(\U1/aes_core/n138 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U206  ( .A(\U1/rkey_next [38]), .B(
        \U1/aes_core/sc2 [6]), .Y(\U1/aes_core/n139 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U205  ( .A0(\U1/aes_core/n138 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n139 ), .Y(
        \U1/dat_next [38]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U204  ( .A(\U1/rkey_next [39]), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/n136 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U203  ( .A(\U1/rkey_next [39]), .B(
        \U1/aes_core/sc2 [7]), .Y(\U1/aes_core/n137 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U202  ( .A0(\U1/aes_core/n136 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n137 ), .Y(
        \U1/dat_next [39]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U201  ( .A(\U1/rkey_next [3]), .B(
        \U1/aes_core/sb2 [3]), .Y(\U1/aes_core/n134 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U200  ( .A(\U1/rkey_next [3]), .B(
        \U1/aes_core/sc3 [3]), .Y(\U1/aes_core/n135 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U199  ( .A0(\U1/aes_core/n134 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n135 ), .Y(
        \U1/dat_next [3]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U198  ( .A(\U1/rkey_next [40]), .B(
        \U1/aes_core/sb0 [8]), .Y(\U1/aes_core/n132 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U197  ( .A(\U1/rkey_next [40]), .B(
        \U1/aes_core/sc2 [8]), .Y(\U1/aes_core/n133 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U196  ( .A0(\U1/aes_core/n132 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n133 ), .Y(
        \U1/dat_next [40]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U195  ( .A(\U1/rkey_next [41]), .B(
        \U1/aes_core/sb0 [9]), .Y(\U1/aes_core/n130 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U194  ( .A(\U1/rkey_next [41]), .B(
        \U1/aes_core/sc2 [9]), .Y(\U1/aes_core/n131 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U193  ( .A0(\U1/aes_core/n130 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n131 ), .Y(
        \U1/dat_next [41]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U192  ( .A(\U1/rkey_next [42]), .B(
        \U1/aes_core/sb0 [10]), .Y(\U1/aes_core/n128 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U191  ( .A(\U1/rkey_next [42]), .B(
        \U1/aes_core/sc2 [10]), .Y(\U1/aes_core/n129 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U190  ( .A0(\U1/aes_core/n128 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n129 ), .Y(
        \U1/dat_next [42]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U189  ( .A(\U1/rkey_next [43]), .B(
        \U1/aes_core/sb0 [11]), .Y(\U1/aes_core/n126 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U188  ( .A(\U1/rkey_next [43]), .B(
        \U1/aes_core/sc2 [11]), .Y(\U1/aes_core/n127 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U187  ( .A0(\U1/aes_core/n126 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n127 ), .Y(
        \U1/dat_next [43]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U186  ( .A(\U1/rkey_next [44]), .B(
        \U1/aes_core/sb0 [12]), .Y(\U1/aes_core/n124 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U185  ( .A(\U1/rkey_next [44]), .B(
        \U1/aes_core/sc2 [12]), .Y(\U1/aes_core/n125 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U184  ( .A0(\U1/aes_core/n124 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n125 ), .Y(
        \U1/dat_next [44]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U183  ( .A(\U1/rkey_next [45]), .B(
        \U1/aes_core/sb0 [13]), .Y(\U1/aes_core/n122 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U182  ( .A(\U1/rkey_next [45]), .B(
        \U1/aes_core/sc2 [13]), .Y(\U1/aes_core/n123 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U181  ( .A0(\U1/aes_core/n122 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n123 ), .Y(
        \U1/dat_next [45]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U180  ( .A(\U1/rkey_next [46]), .B(
        \U1/aes_core/sb0 [14]), .Y(\U1/aes_core/n120 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U179  ( .A(\U1/rkey_next [46]), .B(
        \U1/aes_core/sc2 [14]), .Y(\U1/aes_core/n121 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U178  ( .A0(\U1/aes_core/n120 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n121 ), .Y(
        \U1/dat_next [46]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U177  ( .A(\U1/rkey_next [47]), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/n118 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U176  ( .A(\U1/rkey_next [47]), .B(
        \U1/aes_core/sc2 [15]), .Y(\U1/aes_core/n119 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U175  ( .A0(\U1/aes_core/n118 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n119 ), .Y(
        \U1/dat_next [47]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U174  ( .A(\U1/rkey_next [48]), .B(
        \U1/aes_core/sb3 [16]), .Y(\U1/aes_core/n116 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U173  ( .A(\U1/rkey_next [48]), .B(
        \U1/aes_core/sc2 [16]), .Y(\U1/aes_core/n117 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U172  ( .A0(\U1/aes_core/n116 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n117 ), .Y(
        \U1/dat_next [48]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U171  ( .A(\U1/rkey_next [49]), .B(
        \U1/aes_core/sb3 [17]), .Y(\U1/aes_core/n114 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U170  ( .A(\U1/rkey_next [49]), .B(
        \U1/aes_core/sc2 [17]), .Y(\U1/aes_core/n115 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U169  ( .A0(\U1/aes_core/n114 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n115 ), .Y(
        \U1/dat_next [49]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U168  ( .A(\U1/rkey_next [4]), .B(
        \U1/aes_core/sb2 [4]), .Y(\U1/aes_core/n112 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U167  ( .A(\U1/rkey_next [4]), .B(
        \U1/aes_core/sc3 [4]), .Y(\U1/aes_core/n113 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U166  ( .A0(\U1/aes_core/n112 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n113 ), .Y(
        \U1/dat_next [4]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U165  ( .A(\U1/rkey_next [50]), .B(
        \U1/aes_core/sb3 [18]), .Y(\U1/aes_core/n110 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U164  ( .A(\U1/rkey_next [50]), .B(
        \U1/aes_core/sc2 [18]), .Y(\U1/aes_core/n111 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U163  ( .A0(\U1/aes_core/n110 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n111 ), .Y(
        \U1/dat_next [50]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U162  ( .A(\U1/rkey_next [51]), .B(
        \U1/aes_core/sb3 [19]), .Y(\U1/aes_core/n108 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U161  ( .A(\U1/rkey_next [51]), .B(
        \U1/aes_core/sc2 [19]), .Y(\U1/aes_core/n109 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U160  ( .A0(\U1/aes_core/n108 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n109 ), .Y(
        \U1/dat_next [51]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U159  ( .A(\U1/rkey_next [52]), .B(
        \U1/aes_core/sb3 [20]), .Y(\U1/aes_core/n106 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U158  ( .A(\U1/rkey_next [52]), .B(
        \U1/aes_core/sc2 [20]), .Y(\U1/aes_core/n107 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U157  ( .A0(\U1/aes_core/n106 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n107 ), .Y(
        \U1/dat_next [52]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U156  ( .A(\U1/rkey_next [53]), .B(
        \U1/aes_core/sb3 [21]), .Y(\U1/aes_core/n104 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U155  ( .A(\U1/rkey_next [53]), .B(
        \U1/aes_core/sc2 [21]), .Y(\U1/aes_core/n105 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U154  ( .A0(\U1/aes_core/n104 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n105 ), .Y(
        \U1/dat_next [53]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U153  ( .A(\U1/rkey_next [54]), .B(
        \U1/aes_core/sb3 [22]), .Y(\U1/aes_core/n102 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U152  ( .A(\U1/rkey_next [54]), .B(
        \U1/aes_core/sc2 [22]), .Y(\U1/aes_core/n103 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U151  ( .A0(\U1/aes_core/n102 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n103 ), .Y(
        \U1/dat_next [54]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U150  ( .A(\U1/rkey_next [55]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/n100 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U149  ( .A(\U1/rkey_next [55]), .B(
        \U1/aes_core/sc2 [23]), .Y(\U1/aes_core/n101 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U148  ( .A0(\U1/aes_core/n100 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n101 ), .Y(
        \U1/dat_next [55]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U147  ( .A(\U1/rkey_next [56]), .B(
        \U1/aes_core/sb2 [24]), .Y(\U1/aes_core/n98 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U146  ( .A(\U1/rkey_next [56]), .B(
        \U1/aes_core/sc2 [24]), .Y(\U1/aes_core/n99 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U145  ( .A0(\U1/aes_core/n98 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n99 ), .Y(
        \U1/dat_next [56]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U144  ( .A(\U1/rkey_next [57]), .B(
        \U1/aes_core/sb2 [25]), .Y(\U1/aes_core/n96 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U143  ( .A(\U1/rkey_next [57]), .B(
        \U1/aes_core/sc2 [25]), .Y(\U1/aes_core/n97 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U142  ( .A0(\U1/aes_core/n96 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n97 ), .Y(
        \U1/dat_next [57]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U141  ( .A(\U1/rkey_next [58]), .B(
        \U1/aes_core/sb2 [26]), .Y(\U1/aes_core/n94 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U140  ( .A(\U1/rkey_next [58]), .B(
        \U1/aes_core/sc2 [26]), .Y(\U1/aes_core/n95 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U139  ( .A0(\U1/aes_core/n94 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n95 ), .Y(
        \U1/dat_next [58]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U138  ( .A(\U1/rkey_next [59]), .B(
        \U1/aes_core/sb2 [27]), .Y(\U1/aes_core/n92 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U137  ( .A(\U1/rkey_next [59]), .B(
        \U1/aes_core/sc2 [27]), .Y(\U1/aes_core/n93 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U136  ( .A0(\U1/aes_core/n92 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n93 ), .Y(
        \U1/dat_next [59]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U135  ( .A(\U1/rkey_next [5]), .B(
        \U1/aes_core/sb2 [5]), .Y(\U1/aes_core/n90 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U134  ( .A(\U1/rkey_next [5]), .B(
        \U1/aes_core/sc3 [5]), .Y(\U1/aes_core/n91 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U133  ( .A0(\U1/aes_core/n90 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n91 ), .Y(
        \U1/dat_next [5]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U132  ( .A(\U1/rkey_next [60]), .B(
        \U1/aes_core/sb2 [28]), .Y(\U1/aes_core/n88 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U131  ( .A(\U1/rkey_next [60]), .B(
        \U1/aes_core/sc2 [28]), .Y(\U1/aes_core/n89 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U130  ( .A0(\U1/aes_core/n88 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n89 ), .Y(
        \U1/dat_next [60]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U129  ( .A(\U1/rkey_next [61]), .B(
        \U1/aes_core/sb2 [29]), .Y(\U1/aes_core/n86 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U128  ( .A(\U1/rkey_next [61]), .B(
        \U1/aes_core/sc2 [29]), .Y(\U1/aes_core/n87 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U127  ( .A0(\U1/aes_core/n86 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n87 ), .Y(
        \U1/dat_next [61]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U126  ( .A(\U1/rkey_next [62]), .B(
        \U1/aes_core/sb2 [30]), .Y(\U1/aes_core/n84 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U125  ( .A(\U1/rkey_next [62]), .B(
        \U1/aes_core/sc2 [30]), .Y(\U1/aes_core/n85 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U124  ( .A0(\U1/aes_core/n84 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n85 ), .Y(
        \U1/dat_next [62]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U123  ( .A(\U1/rkey_next [63]), .B(
        \U1/aes_core/sb2 [31]), .Y(\U1/aes_core/n82 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U122  ( .A(\U1/rkey_next [63]), .B(
        \U1/aes_core/sc2 [31]), .Y(\U1/aes_core/n83 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U121  ( .A0(\U1/aes_core/n82 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n83 ), .Y(
        \U1/dat_next [63]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U120  ( .A(\U1/rkey_next [64]), .B(
        \U1/aes_core/sb0 [0]), .Y(\U1/aes_core/n80 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U119  ( .A(\U1/rkey_next [64]), .B(
        \U1/aes_core/sc1 [0]), .Y(\U1/aes_core/n81 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U118  ( .A0(\U1/aes_core/n80 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n81 ), .Y(
        \U1/dat_next [64]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U117  ( .A(\U1/rkey_next [65]), .B(
        \U1/aes_core/sb0 [1]), .Y(\U1/aes_core/n78 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U116  ( .A(\U1/rkey_next [65]), .B(
        \U1/aes_core/sc1 [1]), .Y(\U1/aes_core/n79 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U115  ( .A0(\U1/aes_core/n78 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n79 ), .Y(
        \U1/dat_next [65]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U114  ( .A(\U1/rkey_next [66]), .B(
        \U1/aes_core/sb0 [2]), .Y(\U1/aes_core/n76 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U113  ( .A(\U1/rkey_next [66]), .B(
        \U1/aes_core/sc1 [2]), .Y(\U1/aes_core/n77 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U112  ( .A0(\U1/aes_core/n76 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n77 ), .Y(
        \U1/dat_next [66]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U111  ( .A(\U1/rkey_next [67]), .B(
        \U1/aes_core/sb0 [3]), .Y(\U1/aes_core/n74 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U110  ( .A(\U1/rkey_next [67]), .B(
        \U1/aes_core/sc1 [3]), .Y(\U1/aes_core/n75 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U109  ( .A0(\U1/aes_core/n74 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n75 ), .Y(
        \U1/dat_next [67]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U108  ( .A(\U1/rkey_next [68]), .B(
        \U1/aes_core/sb0 [4]), .Y(\U1/aes_core/n72 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U107  ( .A(\U1/rkey_next [68]), .B(
        \U1/aes_core/sc1 [4]), .Y(\U1/aes_core/n73 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U106  ( .A0(\U1/aes_core/n72 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n73 ), .Y(
        \U1/dat_next [68]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U105  ( .A(\U1/rkey_next [69]), .B(
        \U1/aes_core/sb0 [5]), .Y(\U1/aes_core/n70 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U104  ( .A(\U1/rkey_next [69]), .B(
        \U1/aes_core/sc1 [5]), .Y(\U1/aes_core/n71 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U103  ( .A0(\U1/aes_core/n70 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n71 ), .Y(
        \U1/dat_next [69]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U102  ( .A(\U1/rkey_next [6]), .B(
        \U1/aes_core/sb2 [6]), .Y(\U1/aes_core/n68 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U101  ( .A(\U1/rkey_next [6]), .B(
        \U1/aes_core/sc3 [6]), .Y(\U1/aes_core/n69 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U100  ( .A0(\U1/aes_core/n68 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n69 ), .Y(
        \U1/dat_next [6]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U99  ( .A(\U1/rkey_next [70]), .B(
        \U1/aes_core/sb0 [6]), .Y(\U1/aes_core/n66 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U98  ( .A(\U1/rkey_next [70]), .B(
        \U1/aes_core/sc1 [6]), .Y(\U1/aes_core/n67 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U97  ( .A0(\U1/aes_core/n66 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n67 ), .Y(
        \U1/dat_next [70]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U96  ( .A(\U1/rkey_next [71]), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/n64 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U95  ( .A(\U1/rkey_next [71]), .B(
        \U1/aes_core/sc1 [7]), .Y(\U1/aes_core/n65 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U94  ( .A0(\U1/aes_core/n64 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n65 ), .Y(
        \U1/dat_next [71]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U93  ( .A(\U1/rkey_next [72]), .B(
        \U1/aes_core/sb3 [8]), .Y(\U1/aes_core/n62 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U92  ( .A(\U1/rkey_next [72]), .B(
        \U1/aes_core/sc1 [8]), .Y(\U1/aes_core/n63 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U91  ( .A0(\U1/aes_core/n62 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n63 ), .Y(
        \U1/dat_next [72]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U90  ( .A(\U1/rkey_next [73]), .B(
        \U1/aes_core/sb3 [9]), .Y(\U1/aes_core/n60 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U89  ( .A(\U1/rkey_next [73]), .B(
        \U1/aes_core/sc1 [9]), .Y(\U1/aes_core/n61 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U88  ( .A0(\U1/aes_core/n60 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n61 ), .Y(
        \U1/dat_next [73]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U87  ( .A(\U1/rkey_next [74]), .B(
        \U1/aes_core/sb3 [10]), .Y(\U1/aes_core/n58 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U86  ( .A(\U1/rkey_next [74]), .B(
        \U1/aes_core/sc1 [10]), .Y(\U1/aes_core/n59 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U85  ( .A0(\U1/aes_core/n58 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n59 ), .Y(
        \U1/dat_next [74]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U84  ( .A(\U1/rkey_next [75]), .B(
        \U1/aes_core/sb3 [11]), .Y(\U1/aes_core/n56 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U83  ( .A(\U1/rkey_next [75]), .B(
        \U1/aes_core/sc1 [11]), .Y(\U1/aes_core/n57 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U82  ( .A0(\U1/aes_core/n56 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n57 ), .Y(
        \U1/dat_next [75]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U81  ( .A(\U1/rkey_next [76]), .B(
        \U1/aes_core/sb3 [12]), .Y(\U1/aes_core/n54 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U80  ( .A(\U1/rkey_next [76]), .B(
        \U1/aes_core/sc1 [12]), .Y(\U1/aes_core/n55 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U79  ( .A0(\U1/aes_core/n54 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n55 ), .Y(
        \U1/dat_next [76]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U78  ( .A(\U1/rkey_next [77]), .B(
        \U1/aes_core/sb3 [13]), .Y(\U1/aes_core/n52 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U77  ( .A(\U1/rkey_next [77]), .B(
        \U1/aes_core/sc1 [13]), .Y(\U1/aes_core/n53 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U76  ( .A0(\U1/aes_core/n52 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n53 ), .Y(
        \U1/dat_next [77]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U75  ( .A(\U1/rkey_next [78]), .B(
        \U1/aes_core/sb3 [14]), .Y(\U1/aes_core/n50 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U74  ( .A(\U1/rkey_next [78]), .B(
        \U1/aes_core/sc1 [14]), .Y(\U1/aes_core/n51 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U73  ( .A0(\U1/aes_core/n50 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n51 ), .Y(
        \U1/dat_next [78]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U72  ( .A(\U1/rkey_next [79]), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/n48 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U71  ( .A(\U1/rkey_next [79]), .B(
        \U1/aes_core/sc1 [15]), .Y(\U1/aes_core/n49 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U70  ( .A0(\U1/aes_core/n48 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n49 ), .Y(
        \U1/dat_next [79]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U69  ( .A(\U1/rkey_next [7]), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/n46 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U68  ( .A(\U1/rkey_next [7]), .B(
        \U1/aes_core/sc3 [7]), .Y(\U1/aes_core/n47 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U67  ( .A0(\U1/aes_core/n46 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n47 ), .Y(
        \U1/dat_next [7]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U66  ( .A(\U1/rkey_next [80]), .B(
        \U1/aes_core/sb2 [16]), .Y(\U1/aes_core/n44 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U65  ( .A(\U1/rkey_next [80]), .B(
        \U1/aes_core/sc1 [16]), .Y(\U1/aes_core/n45 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U64  ( .A0(\U1/aes_core/n44 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n45 ), .Y(
        \U1/dat_next [80]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U63  ( .A(\U1/rkey_next [81]), .B(
        \U1/aes_core/sb2 [17]), .Y(\U1/aes_core/n42 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U62  ( .A(\U1/rkey_next [81]), .B(
        \U1/aes_core/sc1 [17]), .Y(\U1/aes_core/n43 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U61  ( .A0(\U1/aes_core/n42 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n43 ), .Y(
        \U1/dat_next [81]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U60  ( .A(\U1/rkey_next [82]), .B(
        \U1/aes_core/sb2 [18]), .Y(\U1/aes_core/n40 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U59  ( .A(\U1/rkey_next [82]), .B(
        \U1/aes_core/sc1 [18]), .Y(\U1/aes_core/n41 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U58  ( .A0(\U1/aes_core/n40 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n41 ), .Y(
        \U1/dat_next [82]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U57  ( .A(\U1/rkey_next [83]), .B(
        \U1/aes_core/sb2 [19]), .Y(\U1/aes_core/n38 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U56  ( .A(\U1/rkey_next [83]), .B(
        \U1/aes_core/sc1 [19]), .Y(\U1/aes_core/n39 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U55  ( .A0(\U1/aes_core/n38 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n39 ), .Y(
        \U1/dat_next [83]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U54  ( .A(\U1/rkey_next [84]), .B(
        \U1/aes_core/sb2 [20]), .Y(\U1/aes_core/n36 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U53  ( .A(\U1/rkey_next [84]), .B(
        \U1/aes_core/sc1 [20]), .Y(\U1/aes_core/n37 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U52  ( .A0(\U1/aes_core/n36 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n37 ), .Y(
        \U1/dat_next [84]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U51  ( .A(\U1/rkey_next [85]), .B(
        \U1/aes_core/sb2 [21]), .Y(\U1/aes_core/n34 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U50  ( .A(\U1/rkey_next [85]), .B(
        \U1/aes_core/sc1 [21]), .Y(\U1/aes_core/n35 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U49  ( .A0(\U1/aes_core/n34 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n35 ), .Y(
        \U1/dat_next [85]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U48  ( .A(\U1/rkey_next [86]), .B(
        \U1/aes_core/sb2 [22]), .Y(\U1/aes_core/n32 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U47  ( .A(\U1/rkey_next [86]), .B(
        \U1/aes_core/sc1 [22]), .Y(\U1/aes_core/n33 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U46  ( .A0(\U1/aes_core/n32 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n33 ), .Y(
        \U1/dat_next [86]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U45  ( .A(\U1/rkey_next [87]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/n30 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U44  ( .A(\U1/rkey_next [87]), .B(
        \U1/aes_core/sc1 [23]), .Y(\U1/aes_core/n31 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U43  ( .A0(\U1/aes_core/n30 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n31 ), .Y(
        \U1/dat_next [87]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U42  ( .A(\U1/rkey_next [88]), .B(
        \U1/aes_core/sb1 [24]), .Y(\U1/aes_core/n28 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U41  ( .A(\U1/rkey_next [88]), .B(
        \U1/aes_core/sc1 [24]), .Y(\U1/aes_core/n29 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U40  ( .A0(\U1/aes_core/n28 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n29 ), .Y(
        \U1/dat_next [88]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U39  ( .A(\U1/rkey_next [89]), .B(
        \U1/aes_core/sb1 [25]), .Y(\U1/aes_core/n26 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U38  ( .A(\U1/rkey_next [89]), .B(
        \U1/aes_core/sc1 [25]), .Y(\U1/aes_core/n27 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U37  ( .A0(\U1/aes_core/n26 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n27 ), .Y(
        \U1/dat_next [89]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U36  ( .A(\U1/rkey_next [8]), .B(
        \U1/aes_core/sb1 [8]), .Y(\U1/aes_core/n24 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U35  ( .A(\U1/rkey_next [8]), .B(
        \U1/aes_core/sc3 [8]), .Y(\U1/aes_core/n25 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U34  ( .A0(\U1/aes_core/n24 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n25 ), .Y(
        \U1/dat_next [8]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U33  ( .A(\U1/rkey_next [90]), .B(
        \U1/aes_core/sb1 [26]), .Y(\U1/aes_core/n22 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U32  ( .A(\U1/rkey_next [90]), .B(
        \U1/aes_core/sc1 [26]), .Y(\U1/aes_core/n23 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U31  ( .A0(\U1/aes_core/n22 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n23 ), .Y(
        \U1/dat_next [90]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U30  ( .A(\U1/rkey_next [91]), .B(
        \U1/aes_core/sb1 [27]), .Y(\U1/aes_core/n20 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U29  ( .A(\U1/rkey_next [91]), .B(
        \U1/aes_core/sc1 [27]), .Y(\U1/aes_core/n21 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U28  ( .A0(\U1/aes_core/n20 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n21 ), .Y(
        \U1/dat_next [91]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U27  ( .A(\U1/rkey_next [92]), .B(
        \U1/aes_core/sb1 [28]), .Y(\U1/aes_core/n18 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U26  ( .A(\U1/rkey_next [92]), .B(
        \U1/aes_core/sc1 [28]), .Y(\U1/aes_core/n19 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U25  ( .A0(\U1/aes_core/n18 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n19 ), .Y(
        \U1/dat_next [92]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U24  ( .A(\U1/rkey_next [93]), .B(
        \U1/aes_core/sb1 [29]), .Y(\U1/aes_core/n16 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U23  ( .A(\U1/rkey_next [93]), .B(
        \U1/aes_core/sc1 [29]), .Y(\U1/aes_core/n17 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U22  ( .A0(\U1/aes_core/n16 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n17 ), .Y(
        \U1/dat_next [93]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U21  ( .A(\U1/rkey_next [94]), .B(
        \U1/aes_core/sb1 [30]), .Y(\U1/aes_core/n14 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U20  ( .A(\U1/rkey_next [94]), .B(
        \U1/aes_core/sc1 [30]), .Y(\U1/aes_core/n15 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U19  ( .A0(\U1/aes_core/n14 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n15 ), .Y(
        \U1/dat_next [94]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U18  ( .A(\U1/rkey_next [95]), .B(
        \U1/aes_core/sb1 [31]), .Y(\U1/aes_core/n12 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U17  ( .A(\U1/rkey_next [95]), .B(
        \U1/aes_core/sc1 [31]), .Y(\U1/aes_core/n13 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U16  ( .A0(\U1/aes_core/n12 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n13 ), .Y(
        \U1/dat_next [95]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U15  ( .A(\U1/rkey_next [96]), .B(
        \U1/aes_core/sb3 [0]), .Y(\U1/aes_core/n10 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U14  ( .A(\U1/rkey_next [96]), .B(
        \U1/aes_core/sc0 [0]), .Y(\U1/aes_core/n11 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U13  ( .A0(\U1/aes_core/n10 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n11 ), .Y(
        \U1/dat_next [96]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U12  ( .A(\U1/rkey_next [97]), .B(
        \U1/aes_core/sb3 [1]), .Y(\U1/aes_core/n8 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U11  ( .A(\U1/rkey_next [97]), .B(
        \U1/aes_core/sc0 [1]), .Y(\U1/aes_core/n9 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U10  ( .A0(\U1/aes_core/n8 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n9 ), .Y(
        \U1/dat_next [97]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U9  ( .A(\U1/rkey_next [98]), .B(
        \U1/aes_core/sb3 [2]), .Y(\U1/aes_core/n6 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U8  ( .A(\U1/rkey_next [98]), .B(
        \U1/aes_core/sc0 [2]), .Y(\U1/aes_core/n7 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U7  ( .A0(\U1/aes_core/n6 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n7 ), .Y(
        \U1/dat_next [98]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U6  ( .A(\U1/rkey_next [99]), .B(
        \U1/aes_core/sb3 [3]), .Y(\U1/aes_core/n4 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U5  ( .A(\U1/rkey_next [99]), .B(
        \U1/aes_core/sc0 [3]), .Y(\U1/aes_core/n5 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U4  ( .A0(\U1/aes_core/n4 ), .A1(
        \U1/aes_core/n258 ), .B0(\U1/sel ), .B1(\U1/aes_core/n5 ), .Y(
        \U1/dat_next [99]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U3  ( .A(\U1/rkey_next [9]), .B(
        \U1/aes_core/sb1 [9]), .Y(\U1/aes_core/n1 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/U2  ( .A(\U1/rkey_next [9]), .B(
        \U1/aes_core/sc3 [9]), .Y(\U1/aes_core/n3 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/U1  ( .A0(\U1/aes_core/n1 ), .A1(
        \U1/aes_core/n2 ), .B0(\U1/sel ), .B1(\U1/aes_core/n3 ), .Y(
        \U1/dat_next [9]) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U711  ( .A0(\U1/aes_core/SB0/n705 ), .A1(
        \U1/aes_core/SB0/n580 ), .B0(\U1/aes_core/SB0/n582 ), .B1(
        \U1/aes_core/SB0/n597 ), .C0(\U1/aes_core/SB0/n706 ), .Y(
        \U1/aes_core/SB0/n703 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U393  ( .A0(\U1/aes_core/SB0/n209 ), .A1(
        \U1/aes_core/SB0/n1031 ), .B0(\U1/aes_core/SB0/n131 ), .B1(
        \U1/aes_core/SB0/n147 ), .C0(\U1/aes_core/SB0/n361 ), .Y(
        \U1/aes_core/SB0/n1029 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U391  ( .A0(\U1/aes_core/SB0/n1156 ), .A1(
        \U1/aes_core/SB0/n1005 ), .B0(\U1/aes_core/SB0/n1007 ), .B1(
        \U1/aes_core/SB0/n1048 ), .C0(\U1/aes_core/SB0/n1157 ), .Y(
        \U1/aes_core/SB0/n1154 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U363  ( .A0(\U1/aes_core/SB0/n531 ), .A1(
        \U1/aes_core/SB0/n753 ), .B0(\U1/aes_core/SB0/n432 ), .B1(
        \U1/aes_core/SB0/n448 ), .C0(\U1/aes_core/SB0/n683 ), .Y(
        \U1/aes_core/SB0/n751 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U361  ( .A0(\U1/aes_core/SB0/n383 ), .A1(
        \U1/aes_core/SB0/n258 ), .B0(\U1/aes_core/SB0/n260 ), .B1(
        \U1/aes_core/SB0/n275 ), .C0(\U1/aes_core/SB0/n384 ), .Y(
        \U1/aes_core/SB0/n381 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U301  ( .A0(\U1/aes_core/SB0/n956 ), .A1(
        \U1/aes_core/SB0/n1204 ), .B0(\U1/aes_core/SB0/n878 ), .B1(
        \U1/aes_core/SB0/n894 ), .C0(\U1/aes_core/SB0/n1134 ), .Y(
        \U1/aes_core/SB0/n1202 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U300  ( .A0(\U1/aes_core/SB0/n531 ), .A1(
        \U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n432 ), .B1(
        \U1/aes_core/SB0/n434 ), .C0(\U1/aes_core/SB0/n640 ), .Y(
        \U1/aes_core/SB0/n766 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U151  ( .A0(\U1/aes_core/SB0/n209 ), .A1(
        \U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n131 ), .B1(
        \U1/aes_core/SB0/n133 ), .C0(\U1/aes_core/SB0/n318 ), .Y(
        \U1/aes_core/SB0/n1620 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB0/U150  ( .A0(\U1/aes_core/SB0/n956 ), .A1(
        \U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n878 ), .B1(
        \U1/aes_core/SB0/n880 ), .C0(\U1/aes_core/SB0/n1091 ), .Y(
        \U1/aes_core/SB0/n1217 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1724  ( .A(Dout[103]), .B(Dout[102]), .Y(
        \U1/aes_core/SB0/n1672 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1723  ( .A(Dout[101]), .B(Dout[100]), .Y(
        \U1/aes_core/SB0/n1681 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1722  ( .A(\U1/aes_core/SB0/n1672 ), .B(
        \U1/aes_core/SB0/n1681 ), .Y(\U1/aes_core/SB0/n1031 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1721  ( .A(Dout[97]), .Y(
        \U1/aes_core/SB0/n1687 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1720  ( .A(Dout[96]), .Y(
        \U1/aes_core/SB0/n1690 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1719  ( .A(\U1/aes_core/SB0/n1687 ), .B(
        \U1/aes_core/SB0/n1690 ), .Y(\U1/aes_core/SB0/n1680 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1718  ( .A(Dout[99]), .B(Dout[98]), .Y(
        \U1/aes_core/SB0/n1660 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1717  ( .A(\U1/aes_core/SB0/n1680 ), .B(
        \U1/aes_core/SB0/n1660 ), .Y(\U1/aes_core/SB0/n147 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1716  ( .A(\U1/aes_core/SB0/n1031 ), .B(
        \U1/aes_core/SB0/n147 ), .Y(\U1/aes_core/SB0/n340 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U1715  ( .A(Dout[98]), .B(Dout[99]), .Y(
        \U1/aes_core/SB0/n1677 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1714  ( .A(\U1/aes_core/SB0/n1677 ), .B(
        \U1/aes_core/SB0/n1680 ), .Y(\U1/aes_core/SB0/n209 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1713  ( .A(Dout[103]), .Y(
        \U1/aes_core/SB0/n1684 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1712  ( .A(\U1/aes_core/SB0/n1684 ), .B(
        Dout[102]), .Y(\U1/aes_core/SB0/n1654 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1711  ( .A(\U1/aes_core/SB0/n1654 ), .B(
        \U1/aes_core/SB0/n1681 ), .Y(\U1/aes_core/SB0/n1032 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1710  ( .A(\U1/aes_core/SB0/n209 ), .B(
        \U1/aes_core/SB0/n1032 ), .Y(\U1/aes_core/SB0/n243 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1709  ( .A(Dout[99]), .Y(
        \U1/aes_core/SB0/n1689 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U1708  ( .A(Dout[98]), .B(
        \U1/aes_core/SB0/n1689 ), .Y(\U1/aes_core/SB0/n1679 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1707  ( .A(\U1/aes_core/SB0/n1680 ), .B(
        \U1/aes_core/SB0/n1679 ), .Y(\U1/aes_core/SB0/n278 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1706  ( .A(\U1/aes_core/SB0/n278 ), .Y(
        \U1/aes_core/SB0/n113 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1705  ( .A(Dout[100]), .Y(
        \U1/aes_core/SB0/n1688 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1704  ( .A(\U1/aes_core/SB0/n1688 ), .B(
        Dout[101]), .Y(\U1/aes_core/SB0/n1673 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1703  ( .A(Dout[102]), .Y(
        \U1/aes_core/SB0/n1685 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1702  ( .A(\U1/aes_core/SB0/n1685 ), .B(
        Dout[103]), .Y(\U1/aes_core/SB0/n1663 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1701  ( .A(\U1/aes_core/SB0/n1673 ), .B(
        \U1/aes_core/SB0/n1663 ), .Y(\U1/aes_core/SB0/n257 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1700  ( .A(\U1/aes_core/SB0/n257 ), .Y(
        \U1/aes_core/SB0/n159 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1699  ( .A(\U1/aes_core/SB0/n113 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n300 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1698  ( .A(\U1/aes_core/SB0/n1031 ), .Y(
        \U1/aes_core/SB0/n144 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1697  ( .A(Dout[97]), .B(Dout[96]), .Y(
        \U1/aes_core/SB0/n1676 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1696  ( .A(\U1/aes_core/SB0/n1676 ), .B(
        \U1/aes_core/SB0/n1660 ), .Y(\U1/aes_core/SB0/n191 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1695  ( .A(\U1/aes_core/SB0/n191 ), .Y(
        \U1/aes_core/SB0/n103 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1694  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n103 ), .Y(\U1/aes_core/SB0/n186 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1693  ( .A(\U1/aes_core/SB0/n1690 ), .B(
        Dout[97]), .Y(\U1/aes_core/SB0/n1661 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1692  ( .A(\U1/aes_core/SB0/n1679 ), .B(
        \U1/aes_core/SB0/n1661 ), .Y(\U1/aes_core/SB0/n291 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1691  ( .A(\U1/aes_core/SB0/n291 ), .Y(
        \U1/aes_core/SB0/n202 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1690  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n322 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U1689  ( .A(\U1/aes_core/SB0/n300 ), .B(
        \U1/aes_core/SB0/n186 ), .C(\U1/aes_core/SB0/n322 ), .Y(
        \U1/aes_core/SB0/n1641 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1688  ( .A(\U1/aes_core/SB0/n1681 ), .B(
        \U1/aes_core/SB0/n1663 ), .Y(\U1/aes_core/SB0/n258 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1687  ( .A(\U1/aes_core/SB0/n1689 ), .B(
        Dout[98]), .Y(\U1/aes_core/SB0/n1670 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1686  ( .A(\U1/aes_core/SB0/n1670 ), .B(
        \U1/aes_core/SB0/n1661 ), .Y(\U1/aes_core/SB0/n260 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1685  ( .A(\U1/aes_core/SB0/n258 ), .B(
        \U1/aes_core/SB0/n260 ), .Y(\U1/aes_core/SB0/n345 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1684  ( .A(\U1/aes_core/SB0/n1032 ), .Y(
        \U1/aes_core/SB0/n142 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1683  ( .A(Dout[101]), .Y(
        \U1/aes_core/SB0/n1686 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1682  ( .A(\U1/aes_core/SB0/n1688 ), .B(
        \U1/aes_core/SB0/n1686 ), .Y(\U1/aes_core/SB0/n1662 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1681  ( .A(\U1/aes_core/SB0/n1672 ), .B(
        \U1/aes_core/SB0/n1662 ), .Y(\U1/aes_core/SB0/n99 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1680  ( .A(\U1/aes_core/SB0/n99 ), .Y(
        \U1/aes_core/SB0/n168 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1679  ( .A(\U1/aes_core/SB0/n1687 ), .B(
        Dout[96]), .Y(\U1/aes_core/SB0/n1671 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1678  ( .A(\U1/aes_core/SB0/n1671 ), .B(
        \U1/aes_core/SB0/n1660 ), .Y(\U1/aes_core/SB0/n134 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1677  ( .A(\U1/aes_core/SB0/n134 ), .Y(
        \U1/aes_core/SB0/n286 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1676  ( .A0(\U1/aes_core/SB0/n142 ), 
        .A1(\U1/aes_core/SB0/n168 ), .B0(\U1/aes_core/SB0/n286 ), .Y(
        \U1/aes_core/SB0/n1682 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1675  ( .A(\U1/aes_core/SB0/n1676 ), .B(
        \U1/aes_core/SB0/n1679 ), .Y(\U1/aes_core/SB0/n146 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1674  ( .A(\U1/aes_core/SB0/n146 ), .Y(
        \U1/aes_core/SB0/n160 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1673  ( .A(\U1/aes_core/SB0/n1686 ), .B(
        Dout[100]), .Y(\U1/aes_core/SB0/n1655 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1672  ( .A(\U1/aes_core/SB0/n1663 ), .B(
        \U1/aes_core/SB0/n1655 ), .Y(\U1/aes_core/SB0/n106 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1671  ( .A(\U1/aes_core/SB0/n258 ), .B(
        \U1/aes_core/SB0/n106 ), .Y(\U1/aes_core/SB0/n367 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1670  ( .A(\U1/aes_core/SB0/n1684 ), .B(
        \U1/aes_core/SB0/n1685 ), .Y(\U1/aes_core/SB0/n1664 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1669  ( .A(\U1/aes_core/SB0/n1673 ), .B(
        \U1/aes_core/SB0/n1664 ), .Y(\U1/aes_core/SB0/n131 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1668  ( .A(\U1/aes_core/SB0/n131 ), .Y(
        \U1/aes_core/SB0/n387 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1667  ( .A0(\U1/aes_core/SB0/n160 ), 
        .A1(\U1/aes_core/SB0/n367 ), .B0(\U1/aes_core/SB0/n387 ), .B1(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n1683 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1666  ( .AN(\U1/aes_core/SB0/n345 ), 
        .B(\U1/aes_core/SB0/n1682 ), .C(\U1/aes_core/SB0/n1683 ), .Y(
        \U1/aes_core/SB0/n1642 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1665  ( .A(\U1/aes_core/SB0/n1681 ), .B(
        \U1/aes_core/SB0/n1664 ), .Y(\U1/aes_core/SB0/n241 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1664  ( .A(\U1/aes_core/SB0/n1677 ), .B(
        \U1/aes_core/SB0/n1676 ), .Y(\U1/aes_core/SB0/n96 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1663  ( .A(\U1/aes_core/SB0/n1654 ), .B(
        \U1/aes_core/SB0/n1673 ), .Y(\U1/aes_core/SB0/n190 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1662  ( .A(\U1/aes_core/SB0/n1677 ), .B(
        \U1/aes_core/SB0/n1671 ), .Y(\U1/aes_core/SB0/n193 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1661  ( .A(\U1/aes_core/SB0/n1680 ), .B(
        \U1/aes_core/SB0/n1670 ), .Y(\U1/aes_core/SB0/n188 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1660  ( .A(\U1/aes_core/SB0/n188 ), .Y(
        \U1/aes_core/SB0/n208 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1659  ( .A(\U1/aes_core/SB0/n106 ), .Y(
        \U1/aes_core/SB0/n372 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1658  ( .A(\U1/aes_core/SB0/n1679 ), .B(
        \U1/aes_core/SB0/n1671 ), .Y(\U1/aes_core/SB0/n170 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1657  ( .A(\U1/aes_core/SB0/n170 ), .Y(
        \U1/aes_core/SB0/n145 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1656  ( .A0(\U1/aes_core/SB0/n208 ), 
        .A1(\U1/aes_core/SB0/n144 ), .B0(\U1/aes_core/SB0/n372 ), .B1(
        \U1/aes_core/SB0/n145 ), .Y(\U1/aes_core/SB0/n1678 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1655  ( .A0(\U1/aes_core/SB0/n241 ), 
        .A1(\U1/aes_core/SB0/n96 ), .B0(\U1/aes_core/SB0/n190 ), .B1(
        \U1/aes_core/SB0/n193 ), .C0(\U1/aes_core/SB0/n1678 ), .Y(
        \U1/aes_core/SB0/n1643 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1654  ( .A(\U1/aes_core/SB0/n188 ), .B(
        \U1/aes_core/SB0/n241 ), .Y(\U1/aes_core/SB0/n379 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1653  ( .A(\U1/aes_core/SB0/n193 ), .B(
        \U1/aes_core/SB0/n258 ), .Y(\U1/aes_core/SB0/n369 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1652  ( .A(\U1/aes_core/SB0/n369 ), .Y(
        \U1/aes_core/SB0/n1674 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1651  ( .A(\U1/aes_core/SB0/n1677 ), .B(
        \U1/aes_core/SB0/n1661 ), .Y(\U1/aes_core/SB0/n118 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1650  ( .A(\U1/aes_core/SB0/n118 ), .Y(
        \U1/aes_core/SB0/n169 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1649  ( .A(\U1/aes_core/SB0/n1676 ), .B(
        \U1/aes_core/SB0/n1670 ), .Y(\U1/aes_core/SB0/n133 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1648  ( .A(\U1/aes_core/SB0/n133 ), .Y(
        \U1/aes_core/SB0/n122 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1647  ( .A0(\U1/aes_core/SB0/n169 ), 
        .A1(\U1/aes_core/SB0/n122 ), .B0(\U1/aes_core/SB0/n168 ), .Y(
        \U1/aes_core/SB0/n1675 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1646  ( .A(\U1/aes_core/SB0/n1672 ), .B(
        \U1/aes_core/SB0/n1655 ), .Y(\U1/aes_core/SB0/n117 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1645  ( .A(\U1/aes_core/SB0/n117 ), .Y(
        \U1/aes_core/SB0/n167 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1644  ( .A(\U1/aes_core/SB0/n167 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n352 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1643  ( .AN(\U1/aes_core/SB0/n379 ), 
        .B(\U1/aes_core/SB0/n1674 ), .C(\U1/aes_core/SB0/n1675 ), .D(
        \U1/aes_core/SB0/n352 ), .Y(\U1/aes_core/SB0/n1665 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1642  ( .A(\U1/aes_core/SB0/n1662 ), .B(
        \U1/aes_core/SB0/n1664 ), .Y(\U1/aes_core/SB0/n97 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1641  ( .A(\U1/aes_core/SB0/n1672 ), .B(
        \U1/aes_core/SB0/n1673 ), .Y(\U1/aes_core/SB0/n105 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1640  ( .A0(\U1/aes_core/SB0/n1032 ), 
        .A1(\U1/aes_core/SB0/n278 ), .B0(\U1/aes_core/SB0/n97 ), .B1(
        \U1/aes_core/SB0/n188 ), .C0(\U1/aes_core/SB0/n105 ), .C1(
        \U1/aes_core/SB0/n170 ), .Y(\U1/aes_core/SB0/n1666 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1639  ( .A(\U1/aes_core/SB0/n146 ), .B(
        \U1/aes_core/SB0/n1032 ), .Y(\U1/aes_core/SB0/n294 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1638  ( .A(\U1/aes_core/SB0/n372 ), .B(
        \U1/aes_core/SB0/n208 ), .Y(\U1/aes_core/SB0/n341 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1637  ( .A(\U1/aes_core/SB0/n145 ), .B(
        \U1/aes_core/SB0/n144 ), .Y(\U1/aes_core/SB0/n321 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1636  ( .A(\U1/aes_core/SB0/n190 ), .Y(
        \U1/aes_core/SB0/n116 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1635  ( .A(\U1/aes_core/SB0/n116 ), .B(
        \U1/aes_core/SB0/n286 ), .Y(\U1/aes_core/SB0/n283 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1634  ( .AN(\U1/aes_core/SB0/n294 ), 
        .B(\U1/aes_core/SB0/n341 ), .C(\U1/aes_core/SB0/n321 ), .D(
        \U1/aes_core/SB0/n283 ), .Y(\U1/aes_core/SB0/n1667 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1633  ( .A(\U1/aes_core/SB0/n1654 ), .B(
        \U1/aes_core/SB0/n1662 ), .Y(\U1/aes_core/SB0/n371 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1632  ( .A(\U1/aes_core/SB0/n371 ), .B(
        \U1/aes_core/SB0/n134 ), .Y(\U1/aes_core/SB0/n217 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1631  ( .A(\U1/aes_core/SB0/n1670 ), .B(
        \U1/aes_core/SB0/n1671 ), .Y(\U1/aes_core/SB0/n98 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1630  ( .A(\U1/aes_core/SB0/n131 ), .B(
        \U1/aes_core/SB0/n98 ), .Y(\U1/aes_core/SB0/n252 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1629  ( .A(\U1/aes_core/SB0/n252 ), .Y(
        \U1/aes_core/SB0/n1669 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1628  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n286 ), .Y(\U1/aes_core/SB0/n233 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1627  ( .A(\U1/aes_core/SB0/n98 ), .Y(
        \U1/aes_core/SB0/n115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1626  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n115 ), .Y(\U1/aes_core/SB0/n182 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1625  ( .AN(\U1/aes_core/SB0/n217 ), 
        .B(\U1/aes_core/SB0/n1669 ), .C(\U1/aes_core/SB0/n233 ), .D(
        \U1/aes_core/SB0/n182 ), .Y(\U1/aes_core/SB0/n1668 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1624  ( .A(\U1/aes_core/SB0/n1665 ), .B(
        \U1/aes_core/SB0/n1666 ), .C(\U1/aes_core/SB0/n1667 ), .D(
        \U1/aes_core/SB0/n1668 ), .Y(\U1/aes_core/SB0/n450 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1623  ( .A(\U1/aes_core/SB0/n191 ), .B(
        \U1/aes_core/SB0/n371 ), .Y(\U1/aes_core/SB0/n183 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1622  ( .A(\U1/aes_core/SB0/n1655 ), .B(
        \U1/aes_core/SB0/n1664 ), .Y(\U1/aes_core/SB0/n275 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1621  ( .A(\U1/aes_core/SB0/n209 ), .B(
        \U1/aes_core/SB0/n275 ), .Y(\U1/aes_core/SB0/n304 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1620  ( .A(\U1/aes_core/SB0/n97 ), .Y(
        \U1/aes_core/SB0/n141 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1619  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n160 ), .Y(\U1/aes_core/SB0/n355 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1618  ( .A0(\U1/aes_core/SB0/n275 ), 
        .A1(\U1/aes_core/SB0/n98 ), .B0(\U1/aes_core/SB0/n355 ), .Y(
        \U1/aes_core/SB0/n1656 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1617  ( .A(\U1/aes_core/SB0/n260 ), .Y(
        \U1/aes_core/SB0/n165 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1616  ( .A(\U1/aes_core/SB0/n165 ), .B(
        \U1/aes_core/SB0/n142 ), .Y(\U1/aes_core/SB0/n164 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1615  ( .A(\U1/aes_core/SB0/n142 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n205 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1614  ( .A(\U1/aes_core/SB0/n1662 ), .B(
        \U1/aes_core/SB0/n1663 ), .Y(\U1/aes_core/SB0/n135 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1613  ( .A(\U1/aes_core/SB0/n135 ), .Y(
        \U1/aes_core/SB0/n360 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1612  ( .A(\U1/aes_core/SB0/n169 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n336 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1611  ( .A(\U1/aes_core/SB0/n147 ), .Y(
        \U1/aes_core/SB0/n166 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1610  ( .A(\U1/aes_core/SB0/n166 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1609  ( .A(\U1/aes_core/SB0/n164 ), .B(
        \U1/aes_core/SB0/n205 ), .C(\U1/aes_core/SB0/n336 ), .D(
        \U1/aes_core/SB0/n272 ), .Y(\U1/aes_core/SB0/n1657 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1608  ( .A(\U1/aes_core/SB0/n145 ), .B(
        \U1/aes_core/SB0/n167 ), .Y(\U1/aes_core/SB0/n238 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1607  ( .A(\U1/aes_core/SB0/n103 ), .B(
        \U1/aes_core/SB0/n167 ), .Y(\U1/aes_core/SB0/n247 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1606  ( .A(\U1/aes_core/SB0/n105 ), .Y(
        \U1/aes_core/SB0/n112 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1605  ( .A(\U1/aes_core/SB0/n208 ), .B(
        \U1/aes_core/SB0/n112 ), .Y(\U1/aes_core/SB0/n375 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1604  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n169 ), .Y(\U1/aes_core/SB0/n264 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1603  ( .A(\U1/aes_core/SB0/n238 ), .B(
        \U1/aes_core/SB0/n247 ), .C(\U1/aes_core/SB0/n375 ), .D(
        \U1/aes_core/SB0/n264 ), .Y(\U1/aes_core/SB0/n1658 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1602  ( .A(\U1/aes_core/SB0/n193 ), .Y(
        \U1/aes_core/SB0/n224 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1601  ( .A(\U1/aes_core/SB0/n372 ), .B(
        \U1/aes_core/SB0/n224 ), .Y(\U1/aes_core/SB0/n389 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1600  ( .A(\U1/aes_core/SB0/n1660 ), .B(
        \U1/aes_core/SB0/n1661 ), .Y(\U1/aes_core/SB0/n158 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1599  ( .A(\U1/aes_core/SB0/n158 ), .Y(
        \U1/aes_core/SB0/n124 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1598  ( .A(\U1/aes_core/SB0/n372 ), .B(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n324 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1597  ( .A(\U1/aes_core/SB0/n209 ), .Y(
        \U1/aes_core/SB0/n101 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1596  ( .A(\U1/aes_core/SB0/n101 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n289 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1595  ( .A(\U1/aes_core/SB0/n168 ), .B(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n140 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1594  ( .A(\U1/aes_core/SB0/n389 ), .B(
        \U1/aes_core/SB0/n324 ), .C(\U1/aes_core/SB0/n289 ), .D(
        \U1/aes_core/SB0/n140 ), .Y(\U1/aes_core/SB0/n1659 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1593  ( .A(\U1/aes_core/SB0/n183 ), .B(
        \U1/aes_core/SB0/n304 ), .C(\U1/aes_core/SB0/n1656 ), .D(
        \U1/aes_core/SB0/n1657 ), .E(\U1/aes_core/SB0/n1658 ), .F(
        \U1/aes_core/SB0/n1659 ), .Y(\U1/aes_core/SB0/n461 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1592  ( .A(\U1/aes_core/SB0/n461 ), .Y(
        \U1/aes_core/SB0/n1645 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1591  ( .A(\U1/aes_core/SB0/n133 ), .B(
        \U1/aes_core/SB0/n275 ), .Y(\U1/aes_core/SB0/n378 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1590  ( .A(\U1/aes_core/SB0/n1654 ), .B(
        \U1/aes_core/SB0/n1655 ), .Y(\U1/aes_core/SB0/n136 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1589  ( .A(\U1/aes_core/SB0/n136 ), .B(
        \U1/aes_core/SB0/n260 ), .Y(\U1/aes_core/SB0/n251 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1588  ( .A(\U1/aes_core/SB0/n251 ), .Y(
        \U1/aes_core/SB0/n1652 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1587  ( .A(\U1/aes_core/SB0/n258 ), .Y(
        \U1/aes_core/SB0/n111 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1586  ( .A0(\U1/aes_core/SB0/n360 ), 
        .A1(\U1/aes_core/SB0/n111 ), .B0(\U1/aes_core/SB0/n124 ), .Y(
        \U1/aes_core/SB0/n1653 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1585  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n224 ), .Y(\U1/aes_core/SB0/n353 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1584  ( .AN(\U1/aes_core/SB0/n378 ), 
        .B(\U1/aes_core/SB0/n1652 ), .C(\U1/aes_core/SB0/n1653 ), .D(
        \U1/aes_core/SB0/n353 ), .Y(\U1/aes_core/SB0/n1648 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1583  ( .A0(\U1/aes_core/SB0/n147 ), 
        .A1(\U1/aes_core/SB0/n99 ), .B0(\U1/aes_core/SB0/n241 ), .B1(
        \U1/aes_core/SB0/n193 ), .C0(\U1/aes_core/SB0/n134 ), .C1(
        \U1/aes_core/SB0/n117 ), .Y(\U1/aes_core/SB0/n1649 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1582  ( .A(\U1/aes_core/SB0/n99 ), .B(
        \U1/aes_core/SB0/n96 ), .Y(\U1/aes_core/SB0/n313 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1581  ( .A(\U1/aes_core/SB0/n111 ), .B(
        \U1/aes_core/SB0/n169 ), .Y(\U1/aes_core/SB0/n180 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1580  ( .A(\U1/aes_core/SB0/n208 ), .B(
        \U1/aes_core/SB0/n111 ), .Y(\U1/aes_core/SB0/n246 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1579  ( .A(\U1/aes_core/SB0/n224 ), .B(
        \U1/aes_core/SB0/n144 ), .Y(\U1/aes_core/SB0/n374 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1578  ( .AN(\U1/aes_core/SB0/n313 ), 
        .B(\U1/aes_core/SB0/n180 ), .C(\U1/aes_core/SB0/n246 ), .D(
        \U1/aes_core/SB0/n374 ), .Y(\U1/aes_core/SB0/n1650 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1577  ( .A(\U1/aes_core/SB0/n101 ), .B(
        \U1/aes_core/SB0/n116 ), .Y(\U1/aes_core/SB0/n301 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1576  ( .A(\U1/aes_core/SB0/n224 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n234 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1575  ( .A(\U1/aes_core/SB0/n372 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n333 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1574  ( .A(\U1/aes_core/SB0/n165 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n288 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1573  ( .A(\U1/aes_core/SB0/n301 ), .B(
        \U1/aes_core/SB0/n234 ), .C(\U1/aes_core/SB0/n333 ), .D(
        \U1/aes_core/SB0/n288 ), .Y(\U1/aes_core/SB0/n1651 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1572  ( .A(\U1/aes_core/SB0/n1648 ), .B(
        \U1/aes_core/SB0/n1649 ), .C(\U1/aes_core/SB0/n1650 ), .D(
        \U1/aes_core/SB0/n1651 ), .Y(\U1/aes_core/SB0/n1647 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1571  ( .A(\U1/aes_core/SB0/n1647 ), .Y(
        \U1/aes_core/SB0/n119 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1570  ( .A(\U1/aes_core/SB0/n103 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n1646 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1569  ( .AN(\U1/aes_core/SB0/n450 ), 
        .B(\U1/aes_core/SB0/n1645 ), .C(\U1/aes_core/SB0/n119 ), .D(
        \U1/aes_core/SB0/n1646 ), .Y(\U1/aes_core/SB0/n1644 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1568  ( .A(\U1/aes_core/SB0/n340 ), .B(
        \U1/aes_core/SB0/n243 ), .C(\U1/aes_core/SB0/n1641 ), .D(
        \U1/aes_core/SB0/n1642 ), .E(\U1/aes_core/SB0/n1643 ), .F(
        \U1/aes_core/SB0/n1644 ), .Y(\U1/aes_core/SB0/n1012 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1567  ( .A(\U1/aes_core/SB0/n118 ), .B(
        \U1/aes_core/SB0/n1032 ), .Y(\U1/aes_core/SB0/n295 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1566  ( .A(\U1/aes_core/SB0/n168 ), .B(
        \U1/aes_core/SB0/n101 ), .Y(\U1/aes_core/SB0/n244 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1565  ( .A(\U1/aes_core/SB0/n112 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n342 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1564  ( .A(\U1/aes_core/SB0/n371 ), .Y(
        \U1/aes_core/SB0/n123 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1563  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n319 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1562  ( .AN(\U1/aes_core/SB0/n295 ), 
        .B(\U1/aes_core/SB0/n244 ), .C(\U1/aes_core/SB0/n342 ), .D(
        \U1/aes_core/SB0/n319 ), .Y(\U1/aes_core/SB0/n1634 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1561  ( .A(\U1/aes_core/SB0/n131 ), .B(
        \U1/aes_core/SB0/n260 ), .Y(\U1/aes_core/SB0/n218 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1560  ( .A(\U1/aes_core/SB0/n208 ), .B(
        \U1/aes_core/SB0/n142 ), .Y(\U1/aes_core/SB0/n362 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1559  ( .A0(\U1/aes_core/SB0/n122 ), 
        .A1(\U1/aes_core/SB0/n202 ), .B0(\U1/aes_core/SB0/n372 ), .Y(
        \U1/aes_core/SB0/n1640 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1558  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n270 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1557  ( .AN(\U1/aes_core/SB0/n218 ), 
        .B(\U1/aes_core/SB0/n362 ), .C(\U1/aes_core/SB0/n1640 ), .D(
        \U1/aes_core/SB0/n270 ), .Y(\U1/aes_core/SB0/n1639 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1556  ( .A(\U1/aes_core/SB0/n1639 ), .Y(
        \U1/aes_core/SB0/n1635 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1555  ( .A(\U1/aes_core/SB0/n241 ), .Y(
        \U1/aes_core/SB0/n121 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1554  ( .A(\U1/aes_core/SB0/n96 ), .Y(
        \U1/aes_core/SB0/n201 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U1553  ( .A0(\U1/aes_core/SB0/n101 ), 
        .A1(\U1/aes_core/SB0/n167 ), .B0(\U1/aes_core/SB0/n121 ), .B1(
        \U1/aes_core/SB0/n286 ), .C0(\U1/aes_core/SB0/n201 ), .C1(
        \U1/aes_core/SB0/n123 ), .Y(\U1/aes_core/SB0/n1636 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1552  ( .A0(\U1/aes_core/SB0/n275 ), 
        .A1(\U1/aes_core/SB0/n118 ), .B0(\U1/aes_core/SB0/n98 ), .B1(
        \U1/aes_core/SB0/n97 ), .Y(\U1/aes_core/SB0/n1638 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1551  ( .A0(\U1/aes_core/SB0/n224 ), 
        .A1(\U1/aes_core/SB0/n387 ), .B0(\U1/aes_core/SB0/n168 ), .B1(
        \U1/aes_core/SB0/n145 ), .C0(\U1/aes_core/SB0/n1638 ), .Y(
        \U1/aes_core/SB0/n1637 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1550  ( .AN(\U1/aes_core/SB0/n1634 ), 
        .B(\U1/aes_core/SB0/n1635 ), .C(\U1/aes_core/SB0/n1636 ), .D(
        \U1/aes_core/SB0/n1637 ), .Y(\U1/aes_core/SB0/n452 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1549  ( .A(\U1/aes_core/SB0/n97 ), .B(
        \U1/aes_core/SB0/n260 ), .Y(\U1/aes_core/SB0/n377 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1548  ( .A0(\U1/aes_core/SB0/n190 ), 
        .A1(\U1/aes_core/SB0/n97 ), .B0(\U1/aes_core/SB0/n158 ), .Y(
        \U1/aes_core/SB0/n1629 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1547  ( .A(\U1/aes_core/SB0/n158 ), .B(
        \U1/aes_core/SB0/n170 ), .Y(\U1/aes_core/SB0/n293 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB0/U1546  ( .A0(\U1/aes_core/SB0/n169 ), .A1(
        \U1/aes_core/SB0/n387 ), .B0(\U1/aes_core/SB0/n293 ), .B1(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n1630 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1545  ( .A0(\U1/aes_core/SB0/n136 ), 
        .A1(\U1/aes_core/SB0/n96 ), .B0(\U1/aes_core/SB0/n371 ), .B1(
        \U1/aes_core/SB0/n278 ), .C0(\U1/aes_core/SB0/n134 ), .C1(
        \U1/aes_core/SB0/n105 ), .Y(\U1/aes_core/SB0/n1631 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1544  ( .A(\U1/aes_core/SB0/n275 ), .Y(
        \U1/aes_core/SB0/n207 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1543  ( .A(\U1/aes_core/SB0/n103 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n181 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1542  ( .A(\U1/aes_core/SB0/n208 ), .B(
        \U1/aes_core/SB0/n387 ), .Y(\U1/aes_core/SB0/n354 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1541  ( .A(\U1/aes_core/SB0/n372 ), .B(
        \U1/aes_core/SB0/n165 ), .Y(\U1/aes_core/SB0/n334 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1540  ( .A(\U1/aes_core/SB0/n208 ), .B(
        \U1/aes_core/SB0/n167 ), .Y(\U1/aes_core/SB0/n235 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1539  ( .A(\U1/aes_core/SB0/n181 ), .B(
        \U1/aes_core/SB0/n354 ), .C(\U1/aes_core/SB0/n334 ), .D(
        \U1/aes_core/SB0/n235 ), .Y(\U1/aes_core/SB0/n1632 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1538  ( .A(\U1/aes_core/SB0/n188 ), .B(
        \U1/aes_core/SB0/n275 ), .Y(\U1/aes_core/SB0/n312 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1537  ( .A(\U1/aes_core/SB0/n202 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n302 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1536  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n286 ), .Y(\U1/aes_core/SB0/n271 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1535  ( .AN(\U1/aes_core/SB0/n312 ), 
        .B(\U1/aes_core/SB0/n302 ), .C(\U1/aes_core/SB0/n271 ), .Y(
        \U1/aes_core/SB0/n1633 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1534  ( .A(\U1/aes_core/SB0/n377 ), .B(
        \U1/aes_core/SB0/n1629 ), .C(\U1/aes_core/SB0/n1630 ), .D(
        \U1/aes_core/SB0/n1631 ), .E(\U1/aes_core/SB0/n1632 ), .F(
        \U1/aes_core/SB0/n1633 ), .Y(\U1/aes_core/SB0/n90 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1533  ( .A0(\U1/aes_core/SB0/n372 ), 
        .A1(\U1/aes_core/SB0/n144 ), .B0(\U1/aes_core/SB0/n113 ), .Y(
        \U1/aes_core/SB0/n1628 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1532  ( .A(\U1/aes_core/SB0/n387 ), .B(
        \U1/aes_core/SB0/n286 ), .Y(\U1/aes_core/SB0/n249 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1531  ( .A(\U1/aes_core/SB0/n169 ), .B(
        \U1/aes_core/SB0/n121 ), .Y(\U1/aes_core/SB0/n357 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1530  ( .A(\U1/aes_core/SB0/n121 ), .B(
        \U1/aes_core/SB0/n165 ), .Y(\U1/aes_core/SB0/n306 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1529  ( .A(\U1/aes_core/SB0/n1628 ), .B(
        \U1/aes_core/SB0/n249 ), .C(\U1/aes_core/SB0/n357 ), .D(
        \U1/aes_core/SB0/n306 ), .Y(\U1/aes_core/SB0/n1624 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1528  ( .A0(\U1/aes_core/SB0/n118 ), 
        .A1(\U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n371 ), .B1(
        \U1/aes_core/SB0/n146 ), .C0(\U1/aes_core/SB0/n117 ), .C1(
        \U1/aes_core/SB0/n260 ), .Y(\U1/aes_core/SB0/n1625 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1527  ( .A(\U1/aes_core/SB0/n166 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n325 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1526  ( .A(\U1/aes_core/SB0/n167 ), .B(
        \U1/aes_core/SB0/n115 ), .Y(\U1/aes_core/SB0/n185 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1525  ( .A(\U1/aes_core/SB0/n167 ), .B(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n338 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1524  ( .A(\U1/aes_core/SB0/n112 ), .B(
        \U1/aes_core/SB0/n122 ), .Y(\U1/aes_core/SB0/n376 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1523  ( .A(\U1/aes_core/SB0/n325 ), .B(
        \U1/aes_core/SB0/n185 ), .C(\U1/aes_core/SB0/n338 ), .D(
        \U1/aes_core/SB0/n376 ), .Y(\U1/aes_core/SB0/n1626 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1522  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n263 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1521  ( .A(\U1/aes_core/SB0/n103 ), .B(
        \U1/aes_core/SB0/n142 ), .Y(\U1/aes_core/SB0/n290 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1520  ( .A(\U1/aes_core/SB0/n113 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n239 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1519  ( .A(\U1/aes_core/SB0/n360 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n390 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1518  ( .A(\U1/aes_core/SB0/n263 ), .B(
        \U1/aes_core/SB0/n290 ), .C(\U1/aes_core/SB0/n239 ), .D(
        \U1/aes_core/SB0/n390 ), .Y(\U1/aes_core/SB0/n1627 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1517  ( .A(\U1/aes_core/SB0/n1624 ), .B(
        \U1/aes_core/SB0/n1625 ), .C(\U1/aes_core/SB0/n1626 ), .D(
        \U1/aes_core/SB0/n1627 ), .Y(\U1/aes_core/SB0/n463 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1516  ( .A(\U1/aes_core/SB0/n1012 ), .B(
        \U1/aes_core/SB0/n452 ), .C(\U1/aes_core/SB0/n90 ), .D(
        \U1/aes_core/SB0/n463 ), .Y(\U1/aes_core/SB0/n1614 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1515  ( .A(\U1/aes_core/SB0/n136 ), .Y(
        \U1/aes_core/SB0/n212 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1514  ( .A0(\U1/aes_core/SB0/n260 ), 
        .A1(\U1/aes_core/SB0/n1031 ), .B0(\U1/aes_core/SB0/n291 ), .B1(
        \U1/aes_core/SB0/n105 ), .Y(\U1/aes_core/SB0/n1623 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1513  ( .A0(\U1/aes_core/SB0/n212 ), 
        .A1(\U1/aes_core/SB0/n160 ), .B0(\U1/aes_core/SB0/n111 ), .B1(
        \U1/aes_core/SB0/n103 ), .C0(\U1/aes_core/SB0/n1623 ), .Y(
        \U1/aes_core/SB0/n1615 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1512  ( .A(\U1/aes_core/SB0/n191 ), .B(
        \U1/aes_core/SB0/n188 ), .Y(\U1/aes_core/SB0/n192 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1511  ( .A0(\U1/aes_core/SB0/n257 ), 
        .A1(\U1/aes_core/SB0/n188 ), .B0(\U1/aes_core/SB0/n275 ), .B1(
        \U1/aes_core/SB0/n147 ), .Y(\U1/aes_core/SB0/n1622 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1510  ( .A0(\U1/aes_core/SB0/n360 ), 
        .A1(\U1/aes_core/SB0/n192 ), .B0(\U1/aes_core/SB0/n141 ), .B1(
        \U1/aes_core/SB0/n122 ), .C0(\U1/aes_core/SB0/n1622 ), .Y(
        \U1/aes_core/SB0/n1616 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1509  ( .A(\U1/aes_core/SB0/n117 ), .B(
        \U1/aes_core/SB0/n258 ), .Y(\U1/aes_core/SB0/n1618 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1508  ( .A(\U1/aes_core/SB0/n167 ), .B(
        \U1/aes_core/SB0/n142 ), .Y(\U1/aes_core/SB0/n200 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1507  ( .A(\U1/aes_core/SB0/n200 ), .Y(
        \U1/aes_core/SB0/n1619 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1506  ( .A(\U1/aes_core/SB0/n209 ), .B(
        \U1/aes_core/SB0/n136 ), .Y(\U1/aes_core/SB0/n328 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1505  ( .A(\U1/aes_core/SB0/n131 ), .B(
        \U1/aes_core/SB0/n133 ), .Y(\U1/aes_core/SB0/n175 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1503  ( .A(\U1/aes_core/SB0/n160 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n318 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1501  ( .A0(\U1/aes_core/SB0/n201 ), 
        .A1(\U1/aes_core/SB0/n1618 ), .B0(\U1/aes_core/SB0/n224 ), .B1(
        \U1/aes_core/SB0/n1619 ), .C0(\U1/aes_core/SB0/n1620 ), .Y(
        \U1/aes_core/SB0/n1617 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1500  ( .AN(\U1/aes_core/SB0/n1614 ), 
        .B(\U1/aes_core/SB0/n1615 ), .C(\U1/aes_core/SB0/n1616 ), .D(
        \U1/aes_core/SB0/n1617 ), .Y(\U1/aes_core/sb0 [0]) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1499  ( .A(Dout[110]), .Y(
        \U1/aes_core/SB0/n1607 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1498  ( .A(Dout[111]), .Y(
        \U1/aes_core/SB0/n1612 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1497  ( .A(\U1/aes_core/SB0/n1607 ), .B(
        \U1/aes_core/SB0/n1612 ), .Y(\U1/aes_core/SB0/n1602 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1496  ( .A(Dout[109]), .Y(
        \U1/aes_core/SB0/n1613 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1495  ( .A(\U1/aes_core/SB0/n1613 ), .B(
        Dout[108]), .Y(\U1/aes_core/SB0/n1595 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1494  ( .A(\U1/aes_core/SB0/n1602 ), .B(
        \U1/aes_core/SB0/n1595 ), .Y(\U1/aes_core/SB0/n54 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1493  ( .A(Dout[107]), .Y(
        \U1/aes_core/SB0/n1604 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1492  ( .A(\U1/aes_core/SB0/n1604 ), .B(
        Dout[106]), .Y(\U1/aes_core/SB0/n1589 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1491  ( .A(Dout[104]), .Y(
        \U1/aes_core/SB0/n1611 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1490  ( .A(\U1/aes_core/SB0/n1611 ), .B(
        Dout[105]), .Y(\U1/aes_core/SB0/n1601 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1489  ( .A(\U1/aes_core/SB0/n1589 ), .B(
        \U1/aes_core/SB0/n1601 ), .Y(\U1/aes_core/SB0/n1450 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1488  ( .A(\U1/aes_core/SB0/n54 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1541 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1487  ( .A(Dout[105]), .Y(
        \U1/aes_core/SB0/n1610 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1486  ( .A(\U1/aes_core/SB0/n1610 ), .B(
        Dout[104]), .Y(\U1/aes_core/SB0/n1592 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1485  ( .A(Dout[106]), .Y(
        \U1/aes_core/SB0/n1605 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1484  ( .A(\U1/aes_core/SB0/n1605 ), .B(
        Dout[107]), .Y(\U1/aes_core/SB0/n1608 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1483  ( .A(\U1/aes_core/SB0/n1592 ), .B(
        \U1/aes_core/SB0/n1608 ), .Y(\U1/aes_core/SB0/n8 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1482  ( .A(Dout[108]), .Y(
        \U1/aes_core/SB0/n1609 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1481  ( .A(\U1/aes_core/SB0/n1613 ), .B(
        \U1/aes_core/SB0/n1609 ), .Y(\U1/aes_core/SB0/n1581 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1480  ( .A(\U1/aes_core/SB0/n1612 ), .B(
        Dout[110]), .Y(\U1/aes_core/SB0/n1606 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1479  ( .A(\U1/aes_core/SB0/n1581 ), .B(
        \U1/aes_core/SB0/n1606 ), .Y(\U1/aes_core/SB0/n1341 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1478  ( .A0(\U1/aes_core/SB0/n1450 ), 
        .A1(\U1/aes_core/SB0/n8 ), .B0(\U1/aes_core/SB0/n1341 ), .Y(
        \U1/aes_core/SB0/n1596 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1477  ( .A(\U1/aes_core/SB0/n1610 ), .B(
        \U1/aes_core/SB0/n1611 ), .Y(\U1/aes_core/SB0/n1590 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1476  ( .A(\U1/aes_core/SB0/n1608 ), .B(
        \U1/aes_core/SB0/n1590 ), .Y(\U1/aes_core/SB0/n1342 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1475  ( .A(\U1/aes_core/SB0/n1609 ), .B(
        Dout[109]), .Y(\U1/aes_core/SB0/n1579 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1474  ( .A(\U1/aes_core/SB0/n1602 ), .B(
        \U1/aes_core/SB0/n1579 ), .Y(\U1/aes_core/SB0/n1367 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1473  ( .A(Dout[107]), .B(Dout[106]), .Y(
        \U1/aes_core/SB0/n1582 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1472  ( .A(\U1/aes_core/SB0/n1590 ), .B(
        \U1/aes_core/SB0/n1582 ), .Y(\U1/aes_core/SB0/n53 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1471  ( .A(\U1/aes_core/SB0/n53 ), .Y(
        \U1/aes_core/SB0/n15 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1470  ( .A(Dout[105]), .B(Dout[104]), .Y(
        \U1/aes_core/SB0/n1583 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1469  ( .A(\U1/aes_core/SB0/n1608 ), .B(
        \U1/aes_core/SB0/n1583 ), .Y(\U1/aes_core/SB0/n58 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1468  ( .A(\U1/aes_core/SB0/n58 ), .Y(
        \U1/aes_core/SB0/n21 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1467  ( .A(\U1/aes_core/SB0/n15 ), .B(
        \U1/aes_core/SB0/n21 ), .Y(\U1/aes_core/SB0/n1539 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1466  ( .A(Dout[111]), .B(Dout[110]), .Y(
        \U1/aes_core/SB0/n1588 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1465  ( .A(\U1/aes_core/SB0/n1595 ), .B(
        \U1/aes_core/SB0/n1588 ), .Y(\U1/aes_core/SB0/n45 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1464  ( .A0(\U1/aes_core/SB0/n1342 ), 
        .A1(\U1/aes_core/SB0/n1367 ), .B0(\U1/aes_core/SB0/n1539 ), .B1(
        \U1/aes_core/SB0/n45 ), .Y(\U1/aes_core/SB0/n1597 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1463  ( .A(\U1/aes_core/SB0/n1608 ), .B(
        \U1/aes_core/SB0/n1601 ), .Y(\U1/aes_core/SB0/n1474 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1462  ( .A(\U1/aes_core/SB0/n1595 ), .B(
        \U1/aes_core/SB0/n1606 ), .Y(\U1/aes_core/SB0/n10 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1461  ( .A(Dout[109]), .B(Dout[108]), .Y(
        \U1/aes_core/SB0/n1603 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1460  ( .A(\U1/aes_core/SB0/n1602 ), .B(
        \U1/aes_core/SB0/n1603 ), .Y(\U1/aes_core/SB0/n74 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1459  ( .A(\U1/aes_core/SB0/n1579 ), .B(
        \U1/aes_core/SB0/n1606 ), .Y(\U1/aes_core/SB0/n76 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1458  ( .A(\U1/aes_core/SB0/n1589 ), .B(
        \U1/aes_core/SB0/n1583 ), .Y(\U1/aes_core/SB0/n1352 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1457  ( .A0(\U1/aes_core/SB0/n1474 ), 
        .A1(\U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n53 ), .B1(
        \U1/aes_core/SB0/n74 ), .C0(\U1/aes_core/SB0/n76 ), .C1(
        \U1/aes_core/SB0/n1352 ), .Y(\U1/aes_core/SB0/n1598 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1456  ( .A(\U1/aes_core/SB0/n1607 ), .B(
        Dout[111]), .Y(\U1/aes_core/SB0/n1580 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1455  ( .A(\U1/aes_core/SB0/n1580 ), .B(
        \U1/aes_core/SB0/n1603 ), .Y(\U1/aes_core/SB0/n46 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1454  ( .A(\U1/aes_core/SB0/n46 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1489 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1453  ( .A(\U1/aes_core/SB0/n1592 ), .B(
        \U1/aes_core/SB0/n1589 ), .Y(\U1/aes_core/SB0/n12 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1452  ( .A(\U1/aes_core/SB0/n12 ), .Y(
        \U1/aes_core/SB0/n1304 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1451  ( .A(\U1/aes_core/SB0/n1603 ), .B(
        \U1/aes_core/SB0/n1606 ), .Y(\U1/aes_core/SB0/n1556 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1450  ( .A(\U1/aes_core/SB0/n1556 ), .Y(
        \U1/aes_core/SB0/n86 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1449  ( .A(\U1/aes_core/SB0/n1304 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n1506 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1448  ( .A(\U1/aes_core/SB0/n1604 ), .B(
        \U1/aes_core/SB0/n1605 ), .Y(\U1/aes_core/SB0/n1593 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1447  ( .A(\U1/aes_core/SB0/n1590 ), .B(
        \U1/aes_core/SB0/n1593 ), .Y(\U1/aes_core/SB0/n1356 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1446  ( .A(\U1/aes_core/SB0/n1356 ), .Y(
        \U1/aes_core/SB0/n1294 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U1445  ( .A(\U1/aes_core/SB0/n1588 ), .B(
        \U1/aes_core/SB0/n1603 ), .Y(\U1/aes_core/SB0/n55 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1444  ( .A(\U1/aes_core/SB0/n1294 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1434 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1443  ( .A(\U1/aes_core/SB0/n1602 ), .B(
        \U1/aes_core/SB0/n1581 ), .Y(\U1/aes_core/SB0/n7 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1442  ( .A(\U1/aes_core/SB0/n7 ), .Y(
        \U1/aes_core/SB0/n49 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1441  ( .A(\U1/aes_core/SB0/n49 ), .B(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n1409 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1440  ( .AN(\U1/aes_core/SB0/n1489 ), 
        .B(\U1/aes_core/SB0/n1506 ), .C(\U1/aes_core/SB0/n1434 ), .D(
        \U1/aes_core/SB0/n1409 ), .Y(\U1/aes_core/SB0/n1599 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1439  ( .A(\U1/aes_core/SB0/n1367 ), .Y(
        \U1/aes_core/SB0/n85 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1438  ( .A(\U1/aes_core/SB0/n1582 ), .B(
        \U1/aes_core/SB0/n1601 ), .Y(\U1/aes_core/SB0/n1345 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1437  ( .A(\U1/aes_core/SB0/n1345 ), .Y(
        \U1/aes_core/SB0/n1308 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1436  ( .A(\U1/aes_core/SB0/n85 ), .B(
        \U1/aes_core/SB0/n1308 ), .Y(\U1/aes_core/SB0/n1519 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1435  ( .A(\U1/aes_core/SB0/n76 ), .Y(
        \U1/aes_core/SB0/n22 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1434  ( .A(\U1/aes_core/SB0/n1601 ), .B(
        \U1/aes_core/SB0/n1593 ), .Y(\U1/aes_core/SB0/n1305 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1433  ( .A(\U1/aes_core/SB0/n1305 ), .Y(
        \U1/aes_core/SB0/n1343 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1432  ( .A(\U1/aes_core/SB0/n22 ), .B(
        \U1/aes_core/SB0/n1343 ), .Y(\U1/aes_core/SB0/n1483 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1431  ( .A(\U1/aes_core/SB0/n85 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1396 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U1430  ( .A(\U1/aes_core/SB0/n1519 ), .B(
        \U1/aes_core/SB0/n1483 ), .C(\U1/aes_core/SB0/n1396 ), .Y(
        \U1/aes_core/SB0/n1600 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1429  ( .A(\U1/aes_core/SB0/n1541 ), .B(
        \U1/aes_core/SB0/n1596 ), .C(\U1/aes_core/SB0/n1597 ), .D(
        \U1/aes_core/SB0/n1598 ), .E(\U1/aes_core/SB0/n1599 ), .F(
        \U1/aes_core/SB0/n1600 ), .Y(\U1/aes_core/SB0/n1 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1428  ( .A(\U1/aes_core/SB0/n1367 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1418 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1427  ( .A(\U1/aes_core/SB0/n1352 ), .Y(
        \U1/aes_core/SB0/n24 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1426  ( .A(\U1/aes_core/SB0/n1474 ), .Y(
        \U1/aes_core/SB0/n20 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1425  ( .A(\U1/aes_core/SB0/n1595 ), .B(
        \U1/aes_core/SB0/n1580 ), .Y(\U1/aes_core/SB0/n11 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1424  ( .A(\U1/aes_core/SB0/n11 ), .Y(
        \U1/aes_core/SB0/n80 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1423  ( .A0(\U1/aes_core/SB0/n24 ), .A1(
        \U1/aes_core/SB0/n20 ), .B0(\U1/aes_core/SB0/n80 ), .Y(
        \U1/aes_core/SB0/n1594 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1422  ( .A(\U1/aes_core/SB0/n49 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1459 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1421  ( .A(\U1/aes_core/SB0/n1341 ), .Y(
        \U1/aes_core/SB0/n1309 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1420  ( .A(\U1/aes_core/SB0/n15 ), .B(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n1497 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1419  ( .AN(\U1/aes_core/SB0/n1418 ), 
        .B(\U1/aes_core/SB0/n1594 ), .C(\U1/aes_core/SB0/n1459 ), .D(
        \U1/aes_core/SB0/n1497 ), .Y(\U1/aes_core/SB0/n1584 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1418  ( .A(\U1/aes_core/SB0/n45 ), .Y(
        \U1/aes_core/SB0/n1386 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1417  ( .A(\U1/aes_core/SB0/n1592 ), .B(
        \U1/aes_core/SB0/n1582 ), .Y(\U1/aes_core/SB0/n1323 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1416  ( .A(\U1/aes_core/SB0/n1323 ), .Y(
        \U1/aes_core/SB0/n14 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1415  ( .A(\U1/aes_core/SB0/n74 ), .Y(
        \U1/aes_core/SB0/n1307 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1414  ( .A(\U1/aes_core/SB0/n1583 ), .B(
        \U1/aes_core/SB0/n1593 ), .Y(\U1/aes_core/SB0/n73 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1413  ( .A(\U1/aes_core/SB0/n73 ), .Y(
        \U1/aes_core/SB0/n23 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U1412  ( .A0(\U1/aes_core/SB0/n1386 ), 
        .A1(\U1/aes_core/SB0/n1294 ), .B0(\U1/aes_core/SB0/n14 ), .B1(
        \U1/aes_core/SB0/n1307 ), .C0(\U1/aes_core/SB0/n23 ), .C1(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n1585 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1411  ( .A(\U1/aes_core/SB0/n54 ), .Y(
        \U1/aes_core/SB0/n1410 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1410  ( .A(\U1/aes_core/SB0/n1588 ), .B(
        \U1/aes_core/SB0/n1581 ), .Y(\U1/aes_core/SB0/n1292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1409  ( .A(\U1/aes_core/SB0/n1592 ), .B(
        \U1/aes_core/SB0/n1593 ), .Y(\U1/aes_core/SB0/n75 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1408  ( .A0(\U1/aes_core/SB0/n1292 ), 
        .A1(\U1/aes_core/SB0/n8 ), .B0(\U1/aes_core/SB0/n75 ), .B1(
        \U1/aes_core/SB0/n1367 ), .Y(\U1/aes_core/SB0/n1591 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1407  ( .A0(\U1/aes_core/SB0/n1304 ), 
        .A1(\U1/aes_core/SB0/n49 ), .B0(\U1/aes_core/SB0/n1410 ), .B1(
        \U1/aes_core/SB0/n1343 ), .C0(\U1/aes_core/SB0/n1591 ), .Y(
        \U1/aes_core/SB0/n1586 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1406  ( .A(\U1/aes_core/SB0/n86 ), .B(
        \U1/aes_core/SB0/n1343 ), .Y(\U1/aes_core/SB0/n1482 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1405  ( .A(\U1/aes_core/SB0/n1589 ), .B(
        \U1/aes_core/SB0/n1590 ), .Y(\U1/aes_core/SB0/n52 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1404  ( .A(\U1/aes_core/SB0/n52 ), .Y(
        \U1/aes_core/SB0/n78 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1403  ( .A(\U1/aes_core/SB0/n78 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n1517 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1402  ( .A(\U1/aes_core/SB0/n1292 ), .Y(
        \U1/aes_core/SB0/n30 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1401  ( .A(\U1/aes_core/SB0/n30 ), .B(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n1433 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1400  ( .A(\U1/aes_core/SB0/n1579 ), .B(
        \U1/aes_core/SB0/n1588 ), .Y(\U1/aes_core/SB0/n1297 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1399  ( .A(\U1/aes_core/SB0/n1297 ), .Y(
        \U1/aes_core/SB0/n32 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1398  ( .A(\U1/aes_core/SB0/n32 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1510 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB0/U1397  ( .A(\U1/aes_core/SB0/n1482 ), .B(
        \U1/aes_core/SB0/n1517 ), .C(\U1/aes_core/SB0/n1433 ), .D(
        \U1/aes_core/SB0/n1510 ), .Y(\U1/aes_core/SB0/n1587 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1396  ( .AN(\U1/aes_core/SB0/n1584 ), 
        .B(\U1/aes_core/SB0/n1585 ), .C(\U1/aes_core/SB0/n1586 ), .D(
        \U1/aes_core/SB0/n1587 ), .Y(\U1/aes_core/SB0/n59 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1395  ( .A(\U1/aes_core/SB0/n1582 ), .B(
        \U1/aes_core/SB0/n1583 ), .Y(\U1/aes_core/SB0/n57 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1394  ( .A(\U1/aes_core/SB0/n57 ), .B(
        \U1/aes_core/SB0/n1341 ), .Y(\U1/aes_core/SB0/n1397 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1393  ( .A(\U1/aes_core/SB0/n54 ), .B(
        \U1/aes_core/SB0/n1356 ), .Y(\U1/aes_core/SB0/n1484 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1392  ( .A(\U1/aes_core/SB0/n21 ), .B(
        \U1/aes_core/SB0/n49 ), .Y(\U1/aes_core/SB0/n1520 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1391  ( .A0(\U1/aes_core/SB0/n54 ), .A1(
        \U1/aes_core/SB0/n12 ), .B0(\U1/aes_core/SB0/n1520 ), .Y(
        \U1/aes_core/SB0/n1575 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1390  ( .A(\U1/aes_core/SB0/n1450 ), .Y(
        \U1/aes_core/SB0/n29 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1389  ( .A(\U1/aes_core/SB0/n86 ), .B(
        \U1/aes_core/SB0/n29 ), .Y(\U1/aes_core/SB0/n1385 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1388  ( .A(\U1/aes_core/SB0/n86 ), .B(
        \U1/aes_core/SB0/n20 ), .Y(\U1/aes_core/SB0/n1408 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1387  ( .A(\U1/aes_core/SB0/n1580 ), .B(
        \U1/aes_core/SB0/n1581 ), .Y(\U1/aes_core/SB0/n1354 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1386  ( .A(\U1/aes_core/SB0/n1354 ), .Y(
        \U1/aes_core/SB0/n47 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1385  ( .A(\U1/aes_core/SB0/n47 ), .B(
        \U1/aes_core/SB0/n1343 ), .Y(\U1/aes_core/SB0/n1507 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1384  ( .A(\U1/aes_core/SB0/n47 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1460 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1383  ( .A(\U1/aes_core/SB0/n1385 ), .B(
        \U1/aes_core/SB0/n1408 ), .C(\U1/aes_core/SB0/n1507 ), .D(
        \U1/aes_core/SB0/n1460 ), .Y(\U1/aes_core/SB0/n1576 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1382  ( .A(\U1/aes_core/SB0/n8 ), .Y(
        \U1/aes_core/SB0/n79 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1381  ( .A(\U1/aes_core/SB0/n79 ), .B(
        \U1/aes_core/SB0/n1386 ), .Y(\U1/aes_core/SB0/n1435 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1380  ( .A(\U1/aes_core/SB0/n57 ), .Y(
        \U1/aes_core/SB0/n72 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1379  ( .A(\U1/aes_core/SB0/n1386 ), .B(
        \U1/aes_core/SB0/n72 ), .Y(\U1/aes_core/SB0/n1440 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1378  ( .A(\U1/aes_core/SB0/n32 ), .B(
        \U1/aes_core/SB0/n78 ), .Y(\U1/aes_core/SB0/n1532 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1377  ( .A(\U1/aes_core/SB0/n55 ), .B(
        \U1/aes_core/SB0/n1343 ), .Y(\U1/aes_core/SB0/n1453 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1376  ( .A(\U1/aes_core/SB0/n1435 ), .B(
        \U1/aes_core/SB0/n1440 ), .C(\U1/aes_core/SB0/n1532 ), .D(
        \U1/aes_core/SB0/n1453 ), .Y(\U1/aes_core/SB0/n1577 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1375  ( .A(\U1/aes_core/SB0/n75 ), .Y(
        \U1/aes_core/SB0/n31 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1374  ( .A(\U1/aes_core/SB0/n80 ), .B(
        \U1/aes_core/SB0/n31 ), .Y(\U1/aes_core/SB0/n1542 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1373  ( .A(\U1/aes_core/SB0/n1308 ), .B(
        \U1/aes_core/SB0/n80 ), .Y(\U1/aes_core/SB0/n1498 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1372  ( .A(\U1/aes_core/SB0/n1579 ), .B(
        \U1/aes_core/SB0/n1580 ), .Y(\U1/aes_core/SB0/n51 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1371  ( .A(\U1/aes_core/SB0/n51 ), .Y(
        \U1/aes_core/SB0/n25 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1370  ( .A(\U1/aes_core/SB0/n1294 ), .B(
        \U1/aes_core/SB0/n25 ), .Y(\U1/aes_core/SB0/n1472 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1369  ( .A(\U1/aes_core/SB0/n1308 ), .B(
        \U1/aes_core/SB0/n30 ), .Y(\U1/aes_core/SB0/n1372 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1368  ( .A(\U1/aes_core/SB0/n1542 ), .B(
        \U1/aes_core/SB0/n1498 ), .C(\U1/aes_core/SB0/n1472 ), .D(
        \U1/aes_core/SB0/n1372 ), .Y(\U1/aes_core/SB0/n1578 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1367  ( .A(\U1/aes_core/SB0/n1397 ), .B(
        \U1/aes_core/SB0/n1484 ), .C(\U1/aes_core/SB0/n1575 ), .D(
        \U1/aes_core/SB0/n1576 ), .E(\U1/aes_core/SB0/n1577 ), .F(
        \U1/aes_core/SB0/n1578 ), .Y(\U1/aes_core/SB0/n68 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1366  ( .A(\U1/aes_core/SB0/n75 ), .B(
        \U1/aes_core/SB0/n1341 ), .Y(\U1/aes_core/SB0/n1531 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1365  ( .A(\U1/aes_core/SB0/n74 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1382 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1364  ( .A(\U1/aes_core/SB0/n76 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1490 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1363  ( .A(\U1/aes_core/SB0/n76 ), .B(
        \U1/aes_core/SB0/n73 ), .Y(\U1/aes_core/SB0/n1481 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1362  ( .A(\U1/aes_core/SB0/n12 ), .B(
        \U1/aes_core/SB0/n46 ), .Y(\U1/aes_core/SB0/n1443 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1361  ( .A(\U1/aes_core/SB0/n47 ), .B(
        \U1/aes_core/SB0/n29 ), .Y(\U1/aes_core/SB0/n1439 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1360  ( .A(\U1/aes_core/SB0/n1304 ), .B(
        \U1/aes_core/SB0/n25 ), .Y(\U1/aes_core/SB0/n1518 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1359  ( .A(\U1/aes_core/SB0/n23 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1505 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1358  ( .AN(\U1/aes_core/SB0/n1443 ), 
        .B(\U1/aes_core/SB0/n1439 ), .C(\U1/aes_core/SB0/n1518 ), .D(
        \U1/aes_core/SB0/n1505 ), .Y(\U1/aes_core/SB0/n1571 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1357  ( .A(\U1/aes_core/SB0/n54 ), .B(
        \U1/aes_core/SB0/n73 ), .Y(\U1/aes_core/SB0/n1471 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1356  ( .A(\U1/aes_core/SB0/n7 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1395 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1355  ( .A(\U1/aes_core/SB0/n1367 ), .B(
        \U1/aes_core/SB0/n8 ), .Y(\U1/aes_core/SB0/n1432 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1354  ( .A(\U1/aes_core/SB0/n1367 ), .B(
        \U1/aes_core/SB0/n1356 ), .Y(\U1/aes_core/SB0/n1534 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1353  ( .A0(\U1/aes_core/SB0/n73 ), .A1(
        \U1/aes_core/SB0/n1367 ), .B0(\U1/aes_core/SB0/n54 ), .B1(
        \U1/aes_core/SB0/n8 ), .Y(\U1/aes_core/SB0/n1573 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1352  ( .A0(\U1/aes_core/SB0/n1474 ), 
        .A1(\U1/aes_core/SB0/n1292 ), .B0(\U1/aes_core/SB0/n1342 ), .B1(
        \U1/aes_core/SB0/n74 ), .Y(\U1/aes_core/SB0/n1574 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1351  ( .A(\U1/aes_core/SB0/n1471 ), .B(
        \U1/aes_core/SB0/n1395 ), .C(\U1/aes_core/SB0/n1432 ), .D(
        \U1/aes_core/SB0/n1534 ), .E(\U1/aes_core/SB0/n1573 ), .F(
        \U1/aes_core/SB0/n1574 ), .Y(\U1/aes_core/SB0/n1572 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1350  ( .A(\U1/aes_core/SB0/n1531 ), .B(
        \U1/aes_core/SB0/n1382 ), .C(\U1/aes_core/SB0/n1490 ), .D(
        \U1/aes_core/SB0/n1481 ), .E(\U1/aes_core/SB0/n1571 ), .F(
        \U1/aes_core/SB0/n1572 ), .Y(\U1/aes_core/SB0/n33 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U1349  ( .A1N(\U1/aes_core/SB0/n55 ), 
        .A0(\U1/aes_core/SB0/n11 ), .B0(\U1/aes_core/SB0/n1342 ), .Y(
        \U1/aes_core/SB0/n1570 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1348  ( .A(\U1/aes_core/SB0/n1367 ), .B(
        \U1/aes_core/SB0/n1323 ), .Y(\U1/aes_core/SB0/n1419 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1347  ( .A(\U1/aes_core/SB0/n74 ), .B(
        \U1/aes_core/SB0/n1305 ), .Y(\U1/aes_core/SB0/n1512 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1346  ( .A(\U1/aes_core/SB0/n74 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1476 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1345  ( .A(\U1/aes_core/SB0/n1570 ), .B(
        \U1/aes_core/SB0/n1419 ), .C(\U1/aes_core/SB0/n1512 ), .D(
        \U1/aes_core/SB0/n1476 ), .Y(\U1/aes_core/SB0/n1565 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1344  ( .A0(\U1/aes_core/SB0/n1305 ), 
        .A1(\U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n1341 ), .B1(
        \U1/aes_core/SB0/n58 ), .C0(\U1/aes_core/SB0/n1450 ), .C1(
        \U1/aes_core/SB0/n45 ), .Y(\U1/aes_core/SB0/n1566 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1343  ( .A(\U1/aes_core/SB0/n12 ), .B(
        \U1/aes_core/SB0/n45 ), .Y(\U1/aes_core/SB0/n1390 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1342  ( .A(\U1/aes_core/SB0/n1297 ), .B(
        \U1/aes_core/SB0/n1352 ), .Y(\U1/aes_core/SB0/n1529 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1341  ( .A(\U1/aes_core/SB0/n1529 ), .Y(
        \U1/aes_core/SB0/n1569 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1340  ( .A(\U1/aes_core/SB0/n25 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1496 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1339  ( .A(\U1/aes_core/SB0/n1386 ), .B(
        \U1/aes_core/SB0/n1308 ), .Y(\U1/aes_core/SB0/n1509 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1338  ( .AN(\U1/aes_core/SB0/n1390 ), 
        .B(\U1/aes_core/SB0/n1569 ), .C(\U1/aes_core/SB0/n1496 ), .D(
        \U1/aes_core/SB0/n1509 ), .Y(\U1/aes_core/SB0/n1567 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1337  ( .A(\U1/aes_core/SB0/n1474 ), .B(
        \U1/aes_core/SB0/n1341 ), .Y(\U1/aes_core/SB0/n1444 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1336  ( .A(\U1/aes_core/SB0/n1556 ), .B(
        \U1/aes_core/SB0/n57 ), .Y(\U1/aes_core/SB0/n1467 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1335  ( .A(\U1/aes_core/SB0/n1354 ), .B(
        \U1/aes_core/SB0/n1342 ), .Y(\U1/aes_core/SB0/n1427 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1334  ( .A(\U1/aes_core/SB0/n1354 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1535 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1333  ( .A(\U1/aes_core/SB0/n1444 ), .B(
        \U1/aes_core/SB0/n1467 ), .C(\U1/aes_core/SB0/n1427 ), .D(
        \U1/aes_core/SB0/n1535 ), .Y(\U1/aes_core/SB0/n1568 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1332  ( .A(\U1/aes_core/SB0/n1565 ), .B(
        \U1/aes_core/SB0/n1566 ), .C(\U1/aes_core/SB0/n1567 ), .D(
        \U1/aes_core/SB0/n1568 ), .Y(\U1/aes_core/SB0/n61 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1331  ( .A(\U1/aes_core/SB0/n46 ), .Y(
        \U1/aes_core/SB0/n27 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1330  ( .A0(\U1/aes_core/SB0/n24 ), .A1(
        \U1/aes_core/SB0/n86 ), .B0(\U1/aes_core/SB0/n1294 ), .B1(
        \U1/aes_core/SB0/n27 ), .Y(\U1/aes_core/SB0/n1564 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1329  ( .A0(\U1/aes_core/SB0/n57 ), 
        .A1(\U1/aes_core/SB0/n7 ), .B0(\U1/aes_core/SB0/n74 ), .B1(
        \U1/aes_core/SB0/n8 ), .C0(\U1/aes_core/SB0/n1564 ), .Y(
        \U1/aes_core/SB0/n1558 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1328  ( .A(\U1/aes_core/SB0/n51 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1500 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1327  ( .A(\U1/aes_core/SB0/n22 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1488 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1326  ( .A(\U1/aes_core/SB0/n86 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1495 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1325  ( .A(\U1/aes_core/SB0/n24 ), .B(
        \U1/aes_core/SB0/n47 ), .Y(\U1/aes_core/SB0/n1523 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1324  ( .AN(\U1/aes_core/SB0/n1500 ), 
        .B(\U1/aes_core/SB0/n1488 ), .C(\U1/aes_core/SB0/n1495 ), .D(
        \U1/aes_core/SB0/n1523 ), .Y(\U1/aes_core/SB0/n1559 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1323  ( .A(\U1/aes_core/SB0/n73 ), .B(
        \U1/aes_core/SB0/n1305 ), .Y(\U1/aes_core/SB0/n1414 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1322  ( .A0(\U1/aes_core/SB0/n29 ), .A1(
        \U1/aes_core/SB0/n1414 ), .B0(\U1/aes_core/SB0/n32 ), .Y(
        \U1/aes_core/SB0/n1561 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1321  ( .A(\U1/aes_core/SB0/n10 ), .Y(
        \U1/aes_core/SB0/n1413 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1320  ( .A0(\U1/aes_core/SB0/n1304 ), 
        .A1(\U1/aes_core/SB0/n31 ), .B0(\U1/aes_core/SB0/n1413 ), .Y(
        \U1/aes_core/SB0/n1562 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1319  ( .A(\U1/aes_core/SB0/n1342 ), .Y(
        \U1/aes_core/SB0/n1302 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1318  ( .A0(\U1/aes_core/SB0/n1410 ), 
        .A1(\U1/aes_core/SB0/n1386 ), .B0(\U1/aes_core/SB0/n1302 ), .Y(
        \U1/aes_core/SB0/n1563 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1317  ( .A(\U1/aes_core/SB0/n1304 ), .B(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n1437 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1316  ( .A(\U1/aes_core/SB0/n1561 ), .B(
        \U1/aes_core/SB0/n1562 ), .C(\U1/aes_core/SB0/n1563 ), .D(
        \U1/aes_core/SB0/n1437 ), .Y(\U1/aes_core/SB0/n1560 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1315  ( .A(\U1/aes_core/SB0/n68 ), .B(
        \U1/aes_core/SB0/n33 ), .C(\U1/aes_core/SB0/n61 ), .D(
        \U1/aes_core/SB0/n1558 ), .E(\U1/aes_core/SB0/n1559 ), .F(
        \U1/aes_core/SB0/n1560 ), .Y(\U1/aes_core/SB0/n1288 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1314  ( .A0(\U1/aes_core/SB0/n1343 ), 
        .A1(\U1/aes_core/SB0/n24 ), .B0(\U1/aes_core/SB0/n30 ), .Y(
        \U1/aes_core/SB0/n1557 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1313  ( .A(\U1/aes_core/SB0/n85 ), .B(
        \U1/aes_core/SB0/n1304 ), .Y(\U1/aes_core/SB0/n1452 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1312  ( .A(\U1/aes_core/SB0/n1307 ), .B(
        \U1/aes_core/SB0/n78 ), .Y(\U1/aes_core/SB0/n1543 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1311  ( .A(\U1/aes_core/SB0/n14 ), .B(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n1441 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1310  ( .A(\U1/aes_core/SB0/n1557 ), .B(
        \U1/aes_core/SB0/n1452 ), .C(\U1/aes_core/SB0/n1543 ), .D(
        \U1/aes_core/SB0/n1441 ), .Y(\U1/aes_core/SB0/n1552 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1309  ( .A0(\U1/aes_core/SB0/n1342 ), 
        .A1(\U1/aes_core/SB0/n1556 ), .B0(\U1/aes_core/SB0/n52 ), .B1(
        \U1/aes_core/SB0/n7 ), .C0(\U1/aes_core/SB0/n8 ), .C1(
        \U1/aes_core/SB0/n1297 ), .Y(\U1/aes_core/SB0/n1553 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1308  ( .A(\U1/aes_core/SB0/n1386 ), .B(
        \U1/aes_core/SB0/n20 ), .Y(\U1/aes_core/SB0/n1521 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1307  ( .A(\U1/aes_core/SB0/n1304 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1398 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1306  ( .A(\U1/aes_core/SB0/n79 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1499 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1305  ( .A(\U1/aes_core/SB0/n14 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1436 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1304  ( .A(\U1/aes_core/SB0/n1521 ), .B(
        \U1/aes_core/SB0/n1398 ), .C(\U1/aes_core/SB0/n1499 ), .D(
        \U1/aes_core/SB0/n1436 ), .Y(\U1/aes_core/SB0/n1554 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1303  ( .A(\U1/aes_core/SB0/n14 ), .B(
        \U1/aes_core/SB0/n22 ), .Y(\U1/aes_core/SB0/n1473 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1302  ( .A(\U1/aes_core/SB0/n21 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n1486 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1301  ( .A(\U1/aes_core/SB0/n80 ), .B(
        \U1/aes_core/SB0/n78 ), .Y(\U1/aes_core/SB0/n1508 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1300  ( .A(\U1/aes_core/SB0/n31 ), .B(
        \U1/aes_core/SB0/n27 ), .Y(\U1/aes_core/SB0/n1533 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1299  ( .A(\U1/aes_core/SB0/n1473 ), .B(
        \U1/aes_core/SB0/n1486 ), .C(\U1/aes_core/SB0/n1508 ), .D(
        \U1/aes_core/SB0/n1533 ), .Y(\U1/aes_core/SB0/n1555 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1298  ( .A(\U1/aes_core/SB0/n1552 ), .B(
        \U1/aes_core/SB0/n1553 ), .C(\U1/aes_core/SB0/n1554 ), .D(
        \U1/aes_core/SB0/n1555 ), .Y(\U1/aes_core/SB0/n1551 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1297  ( .A(\U1/aes_core/SB0/n1551 ), .Y(
        \U1/aes_core/SB0/n70 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1296  ( .A0(\U1/aes_core/SB0/n46 ), 
        .A1(\U1/aes_core/SB0/n1323 ), .B0(\U1/aes_core/SB0/n57 ), .B1(
        \U1/aes_core/SB0/n1292 ), .C0(\U1/aes_core/SB0/n70 ), .Y(
        \U1/aes_core/SB0/n1544 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1295  ( .A(\U1/aes_core/SB0/n25 ), .B(
        \U1/aes_core/SB0/n80 ), .Y(\U1/aes_core/SB0/n1442 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U1294  ( .A1N(\U1/aes_core/SB0/n1442 ), 
        .A0(\U1/aes_core/SB0/n49 ), .B0(\U1/aes_core/SB0/n1343 ), .Y(
        \U1/aes_core/SB0/n1548 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1293  ( .A(\U1/aes_core/SB0/n1345 ), .B(
        \U1/aes_core/SB0/n8 ), .Y(\U1/aes_core/SB0/n1344 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1292  ( .A0(\U1/aes_core/SB0/n23 ), .A1(
        \U1/aes_core/SB0/n1344 ), .B0(\U1/aes_core/SB0/n86 ), .Y(
        \U1/aes_core/SB0/n1549 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1291  ( .A0(\U1/aes_core/SB0/n1304 ), 
        .A1(\U1/aes_core/SB0/n21 ), .B0(\U1/aes_core/SB0/n1307 ), .Y(
        \U1/aes_core/SB0/n1550 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1290  ( .A(\U1/aes_core/SB0/n1308 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1511 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1289  ( .A(\U1/aes_core/SB0/n1548 ), .B(
        \U1/aes_core/SB0/n1549 ), .C(\U1/aes_core/SB0/n1550 ), .D(
        \U1/aes_core/SB0/n1511 ), .Y(\U1/aes_core/SB0/n1545 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1288  ( .A(\U1/aes_core/SB0/n79 ), .B(
        \U1/aes_core/SB0/n1302 ), .Y(\U1/aes_core/SB0/n1303 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1287  ( .A(\U1/aes_core/SB0/n1309 ), .B(
        \U1/aes_core/SB0/n1386 ), .Y(\U1/aes_core/SB0/n1547 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1286  ( .A0(\U1/aes_core/SB0/n1303 ), 
        .A1(\U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n1547 ), .B1(
        \U1/aes_core/SB0/n1352 ), .C0(\U1/aes_core/SB0/n52 ), .C1(
        \U1/aes_core/SB0/n76 ), .Y(\U1/aes_core/SB0/n1546 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1285  ( .A(\U1/aes_core/SB0/n1 ), .B(
        \U1/aes_core/SB0/n59 ), .C(\U1/aes_core/SB0/n1288 ), .D(
        \U1/aes_core/SB0/n1544 ), .E(\U1/aes_core/SB0/n1545 ), .F(
        \U1/aes_core/SB0/n1546 ), .Y(\U1/aes_core/sb0 [10]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1284  ( .A(\U1/aes_core/SB0/n7 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1328 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1283  ( .A(\U1/aes_core/SB0/n24 ), .B(
        \U1/aes_core/SB0/n1410 ), .Y(\U1/aes_core/SB0/n1326 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1282  ( .AN(\U1/aes_core/SB0/n1541 ), 
        .B(\U1/aes_core/SB0/n1542 ), .C(\U1/aes_core/SB0/n1543 ), .D(
        \U1/aes_core/SB0/n1326 ), .Y(\U1/aes_core/SB0/n1536 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1281  ( .A(\U1/aes_core/SB0/n30 ), .B(
        \U1/aes_core/SB0/n1307 ), .Y(\U1/aes_core/SB0/n1379 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1280  ( .A0(\U1/aes_core/SB0/n85 ), .A1(
        \U1/aes_core/SB0/n86 ), .B0(\U1/aes_core/SB0/n31 ), .Y(
        \U1/aes_core/SB0/n1540 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1279  ( .A(\U1/aes_core/SB0/n14 ), .B(
        \U1/aes_core/SB0/n1410 ), .Y(\U1/aes_core/SB0/n1301 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U1278  ( .A0(\U1/aes_core/SB0/n1379 ), 
        .A1(\U1/aes_core/SB0/n58 ), .B0(\U1/aes_core/SB0/n1540 ), .C0(
        \U1/aes_core/SB0/n1301 ), .Y(\U1/aes_core/SB0/n1537 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1277  ( .A0(\U1/aes_core/SB0/n1342 ), 
        .A1(\U1/aes_core/SB0/n1292 ), .B0(\U1/aes_core/SB0/n1539 ), .B1(
        \U1/aes_core/SB0/n46 ), .C0(\U1/aes_core/SB0/n73 ), .C1(
        \U1/aes_core/SB0/n1297 ), .Y(\U1/aes_core/SB0/n1538 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1276  ( .A(\U1/aes_core/SB0/n1534 ), .B(
        \U1/aes_core/SB0/n1328 ), .C(\U1/aes_core/SB0/n1535 ), .D(
        \U1/aes_core/SB0/n1536 ), .E(\U1/aes_core/SB0/n1537 ), .F(
        \U1/aes_core/SB0/n1538 ), .Y(\U1/aes_core/SB0/n1400 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1275  ( .A(\U1/aes_core/SB0/n31 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1322 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1274  ( .AN(\U1/aes_core/SB0/n1531 ), 
        .B(\U1/aes_core/SB0/n1532 ), .C(\U1/aes_core/SB0/n1533 ), .D(
        \U1/aes_core/SB0/n1322 ), .Y(\U1/aes_core/SB0/n1524 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U1273  ( .A0(\U1/aes_core/SB0/n23 ), 
        .A1(\U1/aes_core/SB0/n27 ), .B0(\U1/aes_core/SB0/n22 ), .B1(
        \U1/aes_core/SB0/n20 ), .C0(\U1/aes_core/SB0/n80 ), .C1(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n1525 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1272  ( .A0(\U1/aes_core/SB0/n53 ), .A1(
        \U1/aes_core/SB0/n74 ), .B0(\U1/aes_core/SB0/n1341 ), .B1(
        \U1/aes_core/SB0/n1342 ), .Y(\U1/aes_core/SB0/n1530 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1271  ( .A0(\U1/aes_core/SB0/n1410 ), 
        .A1(\U1/aes_core/SB0/n31 ), .B0(\U1/aes_core/SB0/n78 ), .B1(
        \U1/aes_core/SB0/n55 ), .C0(\U1/aes_core/SB0/n1530 ), .Y(
        \U1/aes_core/SB0/n1526 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1270  ( .A(\U1/aes_core/SB0/n46 ), .B(
        \U1/aes_core/SB0/n11 ), .Y(\U1/aes_core/SB0/n84 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1269  ( .A(\U1/aes_core/SB0/n10 ), .B(
        \U1/aes_core/SB0/n7 ), .Y(\U1/aes_core/SB0/n1528 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1268  ( .A0(\U1/aes_core/SB0/n14 ), 
        .A1(\U1/aes_core/SB0/n84 ), .B0(\U1/aes_core/SB0/n1304 ), .B1(
        \U1/aes_core/SB0/n1528 ), .C0(\U1/aes_core/SB0/n1529 ), .Y(
        \U1/aes_core/SB0/n1527 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1267  ( .AN(\U1/aes_core/SB0/n1524 ), 
        .B(\U1/aes_core/SB0/n1525 ), .C(\U1/aes_core/SB0/n1526 ), .D(
        \U1/aes_core/SB0/n1527 ), .Y(\U1/aes_core/SB0/n1374 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1266  ( .A(\U1/aes_core/SB0/n1367 ), .B(
        \U1/aes_core/SB0/n52 ), .Y(\U1/aes_core/SB0/n1338 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1265  ( .A0(\U1/aes_core/SB0/n51 ), .A1(
        \U1/aes_core/SB0/n52 ), .B0(\U1/aes_core/SB0/n1523 ), .Y(
        \U1/aes_core/SB0/n1513 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1264  ( .A0(\U1/aes_core/SB0/n1304 ), 
        .A1(\U1/aes_core/SB0/n22 ), .B0(\U1/aes_core/SB0/n79 ), .B1(
        \U1/aes_core/SB0/n47 ), .Y(\U1/aes_core/SB0/n1522 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1263  ( .A0(\U1/aes_core/SB0/n10 ), 
        .A1(\U1/aes_core/SB0/n1323 ), .B0(\U1/aes_core/SB0/n1305 ), .B1(
        \U1/aes_core/SB0/n11 ), .C0(\U1/aes_core/SB0/n1522 ), .Y(
        \U1/aes_core/SB0/n1514 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1262  ( .A(\U1/aes_core/SB0/n1450 ), .B(
        \U1/aes_core/SB0/n46 ), .Y(\U1/aes_core/SB0/n62 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1261  ( .A(\U1/aes_core/SB0/n49 ), .B(
        \U1/aes_core/SB0/n31 ), .Y(\U1/aes_core/SB0/n1325 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1260  ( .AN(\U1/aes_core/SB0/n62 ), .B(
        \U1/aes_core/SB0/n1520 ), .C(\U1/aes_core/SB0/n1521 ), .D(
        \U1/aes_core/SB0/n1325 ), .Y(\U1/aes_core/SB0/n1515 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1259  ( .A(\U1/aes_core/SB0/n74 ), .B(
        \U1/aes_core/SB0/n57 ), .Y(\U1/aes_core/SB0/n1347 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1258  ( .AN(\U1/aes_core/SB0/n1347 ), 
        .B(\U1/aes_core/SB0/n1517 ), .C(\U1/aes_core/SB0/n1518 ), .D(
        \U1/aes_core/SB0/n1519 ), .Y(\U1/aes_core/SB0/n1516 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1257  ( .A(\U1/aes_core/SB0/n1338 ), .B(
        \U1/aes_core/SB0/n1512 ), .C(\U1/aes_core/SB0/n1513 ), .D(
        \U1/aes_core/SB0/n1514 ), .E(\U1/aes_core/SB0/n1515 ), .F(
        \U1/aes_core/SB0/n1516 ), .Y(\U1/aes_core/SB0/n1438 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1256  ( .A(\U1/aes_core/SB0/n1345 ), .B(
        \U1/aes_core/SB0/n54 ), .Y(\U1/aes_core/SB0/n1298 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1255  ( .A0(\U1/aes_core/SB0/n1345 ), 
        .A1(\U1/aes_core/SB0/n74 ), .B0(\U1/aes_core/SB0/n1511 ), .Y(
        \U1/aes_core/SB0/n1501 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1254  ( .A(\U1/aes_core/SB0/n11 ), .B(
        \U1/aes_core/SB0/n1450 ), .Y(\U1/aes_core/SB0/n1339 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1253  ( .A(\U1/aes_core/SB0/n1413 ), .B(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n42 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1252  ( .AN(\U1/aes_core/SB0/n1339 ), 
        .B(\U1/aes_core/SB0/n1509 ), .C(\U1/aes_core/SB0/n1510 ), .D(
        \U1/aes_core/SB0/n42 ), .Y(\U1/aes_core/SB0/n1502 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1251  ( .A(\U1/aes_core/SB0/n80 ), .B(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1317 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1250  ( .A(\U1/aes_core/SB0/n15 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n87 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1249  ( .A(\U1/aes_core/SB0/n1343 ), .B(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n19 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1248  ( .A(\U1/aes_core/SB0/n1508 ), .B(
        \U1/aes_core/SB0/n1317 ), .C(\U1/aes_core/SB0/n87 ), .D(
        \U1/aes_core/SB0/n19 ), .Y(\U1/aes_core/SB0/n1503 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1247  ( .A(\U1/aes_core/SB0/n32 ), .B(
        \U1/aes_core/SB0/n21 ), .Y(\U1/aes_core/SB0/n1357 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1246  ( .A(\U1/aes_core/SB0/n1505 ), .B(
        \U1/aes_core/SB0/n1506 ), .C(\U1/aes_core/SB0/n1357 ), .D(
        \U1/aes_core/SB0/n1507 ), .Y(\U1/aes_core/SB0/n1504 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1245  ( .A(\U1/aes_core/SB0/n1298 ), .B(
        \U1/aes_core/SB0/n1500 ), .C(\U1/aes_core/SB0/n1501 ), .D(
        \U1/aes_core/SB0/n1502 ), .E(\U1/aes_core/SB0/n1503 ), .F(
        \U1/aes_core/SB0/n1504 ), .Y(\U1/aes_core/SB0/n1422 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1244  ( .A(\U1/aes_core/SB0/n52 ), .B(
        \U1/aes_core/SB0/n1341 ), .Y(\U1/aes_core/SB0/n1346 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1243  ( .A(\U1/aes_core/SB0/n30 ), .B(
        \U1/aes_core/SB0/n23 ), .Y(\U1/aes_core/SB0/n1321 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1242  ( .A(\U1/aes_core/SB0/n20 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n89 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1241  ( .A(\U1/aes_core/SB0/n1498 ), .B(
        \U1/aes_core/SB0/n1499 ), .C(\U1/aes_core/SB0/n1321 ), .D(
        \U1/aes_core/SB0/n89 ), .Y(\U1/aes_core/SB0/n1491 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1240  ( .A(\U1/aes_core/SB0/n1410 ), .B(
        \U1/aes_core/SB0/n78 ), .Y(\U1/aes_core/SB0/n1335 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1239  ( .A(\U1/aes_core/SB0/n21 ), .B(
        \U1/aes_core/SB0/n1410 ), .Y(\U1/aes_core/SB0/n43 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1238  ( .A(\U1/aes_core/SB0/n1496 ), .B(
        \U1/aes_core/SB0/n1335 ), .C(\U1/aes_core/SB0/n1497 ), .D(
        \U1/aes_core/SB0/n43 ), .Y(\U1/aes_core/SB0/n1492 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U1237  ( .A(\U1/aes_core/SB0/n1307 ), .B(
        \U1/aes_core/SB0/n25 ), .C(\U1/aes_core/SB0/n1309 ), .Y(
        \U1/aes_core/SB0/n1494 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1236  ( .A0(\U1/aes_core/SB0/n1494 ), 
        .A1(\U1/aes_core/SB0/n1352 ), .B0(\U1/aes_core/SB0/n1342 ), .B1(
        \U1/aes_core/SB0/n7 ), .C0(\U1/aes_core/SB0/n1495 ), .Y(
        \U1/aes_core/SB0/n1493 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1235  ( .A(\U1/aes_core/SB0/n1346 ), .B(
        \U1/aes_core/SB0/n1489 ), .C(\U1/aes_core/SB0/n1490 ), .D(
        \U1/aes_core/SB0/n1491 ), .E(\U1/aes_core/SB0/n1492 ), .F(
        \U1/aes_core/SB0/n1493 ), .Y(\U1/aes_core/SB0/n1389 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1234  ( .A(\U1/aes_core/SB0/n54 ), .B(
        \U1/aes_core/SB0/n1474 ), .Y(\U1/aes_core/SB0/n1334 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1233  ( .A0(\U1/aes_core/SB0/n1342 ), 
        .A1(\U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n1488 ), .Y(
        \U1/aes_core/SB0/n1477 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1232  ( .A0(\U1/aes_core/SB0/n1386 ), 
        .A1(\U1/aes_core/SB0/n1343 ), .B0(\U1/aes_core/SB0/n32 ), .B1(
        \U1/aes_core/SB0/n20 ), .Y(\U1/aes_core/SB0/n1487 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1231  ( .A0(\U1/aes_core/SB0/n46 ), 
        .A1(\U1/aes_core/SB0/n8 ), .B0(\U1/aes_core/SB0/n51 ), .B1(
        \U1/aes_core/SB0/n75 ), .C0(\U1/aes_core/SB0/n1487 ), .Y(
        \U1/aes_core/SB0/n1478 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1230  ( .A(\U1/aes_core/SB0/n51 ), .B(
        \U1/aes_core/SB0/n1342 ), .Y(\U1/aes_core/SB0/n63 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1229  ( .A(\U1/aes_core/SB0/n63 ), .Y(
        \U1/aes_core/SB0/n1485 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1228  ( .A(\U1/aes_core/SB0/n22 ), .B(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n1315 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1227  ( .AN(\U1/aes_core/SB0/n1484 ), 
        .B(\U1/aes_core/SB0/n1485 ), .C(\U1/aes_core/SB0/n1486 ), .D(
        \U1/aes_core/SB0/n1315 ), .Y(\U1/aes_core/SB0/n1479 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1226  ( .A(\U1/aes_core/SB0/n1304 ), .B(
        \U1/aes_core/SB0/n47 ), .Y(\U1/aes_core/SB0/n1359 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1225  ( .AN(\U1/aes_core/SB0/n1481 ), 
        .B(\U1/aes_core/SB0/n1482 ), .C(\U1/aes_core/SB0/n1483 ), .D(
        \U1/aes_core/SB0/n1359 ), .Y(\U1/aes_core/SB0/n1480 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1224  ( .A(\U1/aes_core/SB0/n1334 ), .B(
        \U1/aes_core/SB0/n1476 ), .C(\U1/aes_core/SB0/n1477 ), .D(
        \U1/aes_core/SB0/n1478 ), .E(\U1/aes_core/SB0/n1479 ), .F(
        \U1/aes_core/SB0/n1480 ), .Y(\U1/aes_core/SB0/n1415 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1223  ( .A0(\U1/aes_core/SB0/n1309 ), 
        .A1(\U1/aes_core/SB0/n1344 ), .B0(\U1/aes_core/SB0/n1386 ), .B1(
        \U1/aes_core/SB0/n1302 ), .Y(\U1/aes_core/SB0/n1475 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1222  ( .A0(\U1/aes_core/SB0/n73 ), 
        .A1(\U1/aes_core/SB0/n74 ), .B0(\U1/aes_core/SB0/n1474 ), .B1(
        \U1/aes_core/SB0/n11 ), .C0(\U1/aes_core/SB0/n1475 ), .Y(
        \U1/aes_core/SB0/n1464 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1221  ( .A(\U1/aes_core/SB0/n25 ), .B(
        \U1/aes_core/SB0/n29 ), .Y(\U1/aes_core/SB0/n1318 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1220  ( .AN(\U1/aes_core/SB0/n1471 ), 
        .B(\U1/aes_core/SB0/n1472 ), .C(\U1/aes_core/SB0/n1473 ), .D(
        \U1/aes_core/SB0/n1318 ), .Y(\U1/aes_core/SB0/n1465 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1219  ( .A0(\U1/aes_core/SB0/n72 ), .A1(
        \U1/aes_core/SB0/n14 ), .B0(\U1/aes_core/SB0/n32 ), .Y(
        \U1/aes_core/SB0/n1468 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1218  ( .A(\U1/aes_core/SB0/n10 ), .B(
        \U1/aes_core/SB0/n1367 ), .Y(\U1/aes_core/SB0/n1470 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1217  ( .A0(\U1/aes_core/SB0/n21 ), .A1(
        \U1/aes_core/SB0/n1470 ), .B0(\U1/aes_core/SB0/n25 ), .B1(
        \U1/aes_core/SB0/n1414 ), .Y(\U1/aes_core/SB0/n1469 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1216  ( .AN(\U1/aes_core/SB0/n1467 ), 
        .B(\U1/aes_core/SB0/n1468 ), .C(\U1/aes_core/SB0/n1469 ), .Y(
        \U1/aes_core/SB0/n1466 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1215  ( .A(\U1/aes_core/SB0/n1422 ), .B(
        \U1/aes_core/SB0/n1389 ), .C(\U1/aes_core/SB0/n1415 ), .D(
        \U1/aes_core/SB0/n1464 ), .E(\U1/aes_core/SB0/n1465 ), .F(
        \U1/aes_core/SB0/n1466 ), .Y(\U1/aes_core/SB0/n1363 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1214  ( .A(\U1/aes_core/SB0/n1400 ), .B(
        \U1/aes_core/SB0/n1374 ), .C(\U1/aes_core/SB0/n1438 ), .D(
        \U1/aes_core/SB0/n1363 ), .Y(\U1/aes_core/SB0/n1454 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1213  ( .A(\U1/aes_core/SB0/n21 ), .B(
        \U1/aes_core/SB0/n1294 ), .Y(\U1/aes_core/SB0/n1353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1212  ( .A(\U1/aes_core/SB0/n31 ), .B(
        \U1/aes_core/SB0/n1302 ), .Y(\U1/aes_core/SB0/n1360 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1211  ( .A(\U1/aes_core/SB0/n57 ), .B(
        \U1/aes_core/SB0/n52 ), .Y(\U1/aes_core/SB0/n48 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1210  ( .A0(\U1/aes_core/SB0/n1410 ), 
        .A1(\U1/aes_core/SB0/n79 ), .B0(\U1/aes_core/SB0/n48 ), .B1(
        \U1/aes_core/SB0/n49 ), .Y(\U1/aes_core/SB0/n1463 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1209  ( .A0(\U1/aes_core/SB0/n1341 ), 
        .A1(\U1/aes_core/SB0/n1353 ), .B0(\U1/aes_core/SB0/n76 ), .B1(
        \U1/aes_core/SB0/n1360 ), .C0(\U1/aes_core/SB0/n1463 ), .Y(
        \U1/aes_core/SB0/n1462 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1208  ( .A(\U1/aes_core/SB0/n1462 ), .Y(
        \U1/aes_core/SB0/n1455 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1207  ( .A0(\U1/aes_core/SB0/n53 ), .A1(
        \U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n1342 ), .B1(
        \U1/aes_core/SB0/n1367 ), .Y(\U1/aes_core/SB0/n1461 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1206  ( .A0(\U1/aes_core/SB0/n1308 ), 
        .A1(\U1/aes_core/SB0/n86 ), .B0(\U1/aes_core/SB0/n27 ), .B1(
        \U1/aes_core/SB0/n72 ), .C0(\U1/aes_core/SB0/n1461 ), .Y(
        \U1/aes_core/SB0/n1456 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1205  ( .A0(\U1/aes_core/SB0/n1294 ), 
        .A1(\U1/aes_core/SB0/n31 ), .B0(\U1/aes_core/SB0/n1307 ), .Y(
        \U1/aes_core/SB0/n1458 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1204  ( .A(\U1/aes_core/SB0/n14 ), .B(
        \U1/aes_core/SB0/n49 ), .Y(\U1/aes_core/SB0/n1336 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB0/U1203  ( .A(\U1/aes_core/SB0/n1458 ), .B(
        \U1/aes_core/SB0/n1336 ), .C(\U1/aes_core/SB0/n1459 ), .D(
        \U1/aes_core/SB0/n1460 ), .Y(\U1/aes_core/SB0/n1457 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1202  ( .AN(\U1/aes_core/SB0/n1454 ), 
        .B(\U1/aes_core/SB0/n1455 ), .C(\U1/aes_core/SB0/n1456 ), .D(
        \U1/aes_core/SB0/n1457 ), .Y(\U1/aes_core/sb0 [11]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1201  ( .A0(\U1/aes_core/SB0/n1442 ), 
        .A1(\U1/aes_core/SB0/n1354 ), .B0(\U1/aes_core/SB0/n57 ), .Y(
        \U1/aes_core/SB0/n1445 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1200  ( .A(\U1/aes_core/SB0/n1413 ), .B(
        \U1/aes_core/SB0/n29 ), .Y(\U1/aes_core/SB0/n1327 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U1199  ( .A(\U1/aes_core/SB0/n1452 ), .B(
        \U1/aes_core/SB0/n1327 ), .C(\U1/aes_core/SB0/n1453 ), .Y(
        \U1/aes_core/SB0/n1446 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1198  ( .A(\U1/aes_core/SB0/n1309 ), .B(
        \U1/aes_core/SB0/n32 ), .Y(\U1/aes_core/SB0/n1449 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1197  ( .A(\U1/aes_core/SB0/n49 ), .B(
        \U1/aes_core/SB0/n1410 ), .Y(\U1/aes_core/SB0/n1451 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1196  ( .A0(\U1/aes_core/SB0/n1449 ), 
        .A1(\U1/aes_core/SB0/n1450 ), .B0(\U1/aes_core/SB0/n1451 ), .B1(
        \U1/aes_core/SB0/n1305 ), .C0(\U1/aes_core/SB0/n1356 ), .C1(
        \U1/aes_core/SB0/n1354 ), .Y(\U1/aes_core/SB0/n1447 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1195  ( .A0(\U1/aes_core/SB0/n51 ), 
        .A1(\U1/aes_core/SB0/n1345 ), .B0(\U1/aes_core/SB0/n73 ), .B1(
        \U1/aes_core/SB0/n11 ), .C0(\U1/aes_core/SB0/n46 ), .C1(
        \U1/aes_core/SB0/n1352 ), .Y(\U1/aes_core/SB0/n1448 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1194  ( .A(\U1/aes_core/SB0/n1443 ), .B(
        \U1/aes_core/SB0/n1444 ), .C(\U1/aes_core/SB0/n1445 ), .D(
        \U1/aes_core/SB0/n1446 ), .E(\U1/aes_core/SB0/n1447 ), .F(
        \U1/aes_core/SB0/n1448 ), .Y(\U1/aes_core/SB0/n1362 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1193  ( .A0(\U1/aes_core/SB0/n1442 ), 
        .A1(\U1/aes_core/SB0/n74 ), .B0(\U1/aes_core/SB0/n8 ), .Y(
        \U1/aes_core/SB0/n1416 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB0/U1192  ( .A0(\U1/aes_core/SB0/n58 ), .A1(
        \U1/aes_core/SB0/n75 ), .A2(\U1/aes_core/SB0/n1352 ), .B0(
        \U1/aes_core/SB0/n45 ), .Y(\U1/aes_core/SB0/n1417 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1191  ( .A(\U1/aes_core/SB0/n78 ), .B(
        \U1/aes_core/SB0/n27 ), .Y(\U1/aes_core/SB0/n1320 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1190  ( .A(\U1/aes_core/SB0/n1439 ), .B(
        \U1/aes_core/SB0/n1440 ), .C(\U1/aes_core/SB0/n1441 ), .D(
        \U1/aes_core/SB0/n1320 ), .Y(\U1/aes_core/SB0/n1420 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1189  ( .A(\U1/aes_core/SB0/n1438 ), .Y(
        \U1/aes_core/SB0/n1423 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1188  ( .A(\U1/aes_core/SB0/n45 ), .B(
        \U1/aes_core/SB0/n52 ), .Y(\U1/aes_core/SB0/n1340 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1187  ( .A0(\U1/aes_core/SB0/n1360 ), 
        .A1(\U1/aes_core/SB0/n1297 ), .B0(\U1/aes_core/SB0/n1437 ), .Y(
        \U1/aes_core/SB0/n1428 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1186  ( .A0(\U1/aes_core/SB0/n74 ), 
        .A1(\U1/aes_core/SB0/n12 ), .B0(\U1/aes_core/SB0/n57 ), .B1(
        \U1/aes_core/SB0/n1367 ), .C0(\U1/aes_core/SB0/n73 ), .C1(
        \U1/aes_core/SB0/n45 ), .Y(\U1/aes_core/SB0/n1429 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1185  ( .A(\U1/aes_core/SB0/n47 ), .B(
        \U1/aes_core/SB0/n31 ), .Y(\U1/aes_core/SB0/n1316 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1184  ( .A(\U1/aes_core/SB0/n1294 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n82 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1183  ( .A(\U1/aes_core/SB0/n1435 ), .B(
        \U1/aes_core/SB0/n1436 ), .C(\U1/aes_core/SB0/n1316 ), .D(
        \U1/aes_core/SB0/n82 ), .Y(\U1/aes_core/SB0/n1430 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1182  ( .A(\U1/aes_core/SB0/n21 ), .B(
        \U1/aes_core/SB0/n55 ), .Y(\U1/aes_core/SB0/n1358 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1181  ( .AN(\U1/aes_core/SB0/n1432 ), 
        .B(\U1/aes_core/SB0/n1433 ), .C(\U1/aes_core/SB0/n1434 ), .D(
        \U1/aes_core/SB0/n1358 ), .Y(\U1/aes_core/SB0/n1431 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1180  ( .A(\U1/aes_core/SB0/n1340 ), .B(
        \U1/aes_core/SB0/n1427 ), .C(\U1/aes_core/SB0/n1428 ), .D(
        \U1/aes_core/SB0/n1429 ), .E(\U1/aes_core/SB0/n1430 ), .F(
        \U1/aes_core/SB0/n1431 ), .Y(\U1/aes_core/SB0/n1426 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1179  ( .A(\U1/aes_core/SB0/n1426 ), .Y(
        \U1/aes_core/SB0/n1373 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1178  ( .A0(\U1/aes_core/SB0/n10 ), .A1(
        \U1/aes_core/SB0/n1345 ), .B0(\U1/aes_core/SB0/n73 ), .B1(
        \U1/aes_core/SB0/n7 ), .Y(\U1/aes_core/SB0/n1425 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U1177  ( .A0(\U1/aes_core/SB0/n30 ), 
        .A1(\U1/aes_core/SB0/n31 ), .B0(\U1/aes_core/SB0/n24 ), .B1(
        \U1/aes_core/SB0/n55 ), .C0(\U1/aes_core/SB0/n1425 ), .Y(
        \U1/aes_core/SB0/n1424 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1176  ( .AN(\U1/aes_core/SB0/n1422 ), 
        .B(\U1/aes_core/SB0/n1423 ), .C(\U1/aes_core/SB0/n1373 ), .D(
        \U1/aes_core/SB0/n1424 ), .Y(\U1/aes_core/SB0/n1421 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1175  ( .A(\U1/aes_core/SB0/n1416 ), .B(
        \U1/aes_core/SB0/n1417 ), .C(\U1/aes_core/SB0/n1418 ), .D(
        \U1/aes_core/SB0/n1419 ), .E(\U1/aes_core/SB0/n1420 ), .F(
        \U1/aes_core/SB0/n1421 ), .Y(\U1/aes_core/SB0/n1375 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1174  ( .A(\U1/aes_core/SB0/n1415 ), .Y(
        \U1/aes_core/SB0/n1411 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1173  ( .A0(\U1/aes_core/SB0/n1413 ), 
        .A1(\U1/aes_core/SB0/n1414 ), .B0(\U1/aes_core/SB0/n1410 ), .B1(
        \U1/aes_core/SB0/n15 ), .Y(\U1/aes_core/SB0/n1412 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U1172  ( .A0(\U1/aes_core/SB0/n1356 ), 
        .A1(\U1/aes_core/SB0/n45 ), .B0(\U1/aes_core/SB0/n1411 ), .C0(
        \U1/aes_core/SB0/n1412 ), .Y(\U1/aes_core/SB0/n1401 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1171  ( .A0(\U1/aes_core/SB0/n78 ), .A1(
        \U1/aes_core/SB0/n79 ), .B0(\U1/aes_core/SB0/n22 ), .Y(
        \U1/aes_core/SB0/n1406 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1170  ( .A0(\U1/aes_core/SB0/n1410 ), 
        .A1(\U1/aes_core/SB0/n86 ), .B0(\U1/aes_core/SB0/n1302 ), .Y(
        \U1/aes_core/SB0/n1407 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1169  ( .A(\U1/aes_core/SB0/n1406 ), .B(
        \U1/aes_core/SB0/n1407 ), .C(\U1/aes_core/SB0/n1408 ), .D(
        \U1/aes_core/SB0/n1409 ), .Y(\U1/aes_core/SB0/n1402 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1168  ( .A(\U1/aes_core/SB0/n29 ), .B(
        \U1/aes_core/SB0/n20 ), .Y(\U1/aes_core/SB0/n1404 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1167  ( .A(\U1/aes_core/SB0/n23 ), .B(
        \U1/aes_core/SB0/n21 ), .Y(\U1/aes_core/SB0/n1405 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1166  ( .A(\U1/aes_core/SB0/n1386 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n44 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1165  ( .A0(\U1/aes_core/SB0/n1404 ), 
        .A1(\U1/aes_core/SB0/n1292 ), .B0(\U1/aes_core/SB0/n1405 ), .B1(
        \U1/aes_core/SB0/n1354 ), .C0(\U1/aes_core/SB0/n44 ), .C1(
        \U1/aes_core/SB0/n1323 ), .Y(\U1/aes_core/SB0/n1403 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1164  ( .A(\U1/aes_core/SB0/n1362 ), .B(
        \U1/aes_core/SB0/n1375 ), .C(\U1/aes_core/SB0/n1400 ), .D(
        \U1/aes_core/SB0/n1401 ), .E(\U1/aes_core/SB0/n1402 ), .F(
        \U1/aes_core/SB0/n1403 ), .Y(\U1/aes_core/sb0 [12]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1163  ( .A(\U1/aes_core/SB0/n54 ), .B(
        \U1/aes_core/SB0/n57 ), .Y(\U1/aes_core/SB0/n1337 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U1162  ( .A1N(\U1/aes_core/SB0/n48 ), 
        .A0(\U1/aes_core/SB0/n75 ), .B0(\U1/aes_core/SB0/n10 ), .Y(
        \U1/aes_core/SB0/n1391 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1161  ( .A(\U1/aes_core/SB0/n1309 ), .B(
        \U1/aes_core/SB0/n86 ), .Y(\U1/aes_core/SB0/n1399 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1160  ( .A0(\U1/aes_core/SB0/n1292 ), 
        .A1(\U1/aes_core/SB0/n52 ), .B0(\U1/aes_core/SB0/n1399 ), .B1(
        \U1/aes_core/SB0/n73 ), .C0(\U1/aes_core/SB0/n57 ), .C1(
        \U1/aes_core/SB0/n76 ), .Y(\U1/aes_core/SB0/n1392 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1159  ( .A(\U1/aes_core/SB0/n27 ), .B(
        \U1/aes_core/SB0/n1343 ), .Y(\U1/aes_core/SB0/n1319 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1158  ( .A(\U1/aes_core/SB0/n55 ), .B(
        \U1/aes_core/SB0/n72 ), .Y(\U1/aes_core/SB0/n88 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1157  ( .AN(\U1/aes_core/SB0/n1397 ), 
        .B(\U1/aes_core/SB0/n1398 ), .C(\U1/aes_core/SB0/n1319 ), .D(
        \U1/aes_core/SB0/n88 ), .Y(\U1/aes_core/SB0/n1393 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1156  ( .A(\U1/aes_core/SB0/n85 ), .B(
        \U1/aes_core/SB0/n24 ), .Y(\U1/aes_core/SB0/n41 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1155  ( .AN(\U1/aes_core/SB0/n1395 ), 
        .B(\U1/aes_core/SB0/n1396 ), .C(\U1/aes_core/SB0/n41 ), .Y(
        \U1/aes_core/SB0/n1394 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1154  ( .A(\U1/aes_core/SB0/n1337 ), .B(
        \U1/aes_core/SB0/n1390 ), .C(\U1/aes_core/SB0/n1391 ), .D(
        \U1/aes_core/SB0/n1392 ), .E(\U1/aes_core/SB0/n1393 ), .F(
        \U1/aes_core/SB0/n1394 ), .Y(\U1/aes_core/SB0/n1361 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1153  ( .A(\U1/aes_core/SB0/n1389 ), .Y(
        \U1/aes_core/SB0/n1387 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1152  ( .A0(\U1/aes_core/SB0/n32 ), .A1(
        \U1/aes_core/SB0/n1304 ), .B0(\U1/aes_core/SB0/n1302 ), .B1(
        \U1/aes_core/SB0/n27 ), .Y(\U1/aes_core/SB0/n1388 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U1151  ( .A0(\U1/aes_core/SB0/n10 ), 
        .A1(\U1/aes_core/SB0/n8 ), .B0(\U1/aes_core/SB0/n1387 ), .C0(
        \U1/aes_core/SB0/n1388 ), .Y(\U1/aes_core/SB0/n1376 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1150  ( .A0(\U1/aes_core/SB0/n30 ), .A1(
        \U1/aes_core/SB0/n32 ), .B0(\U1/aes_core/SB0/n1343 ), .Y(
        \U1/aes_core/SB0/n1383 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1149  ( .A0(\U1/aes_core/SB0/n29 ), .A1(
        \U1/aes_core/SB0/n15 ), .B0(\U1/aes_core/SB0/n1386 ), .Y(
        \U1/aes_core/SB0/n1384 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1148  ( .AN(\U1/aes_core/SB0/n1382 ), 
        .B(\U1/aes_core/SB0/n1383 ), .C(\U1/aes_core/SB0/n1384 ), .D(
        \U1/aes_core/SB0/n1385 ), .Y(\U1/aes_core/SB0/n1377 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1147  ( .A0(\U1/aes_core/SB0/n22 ), .A1(
        \U1/aes_core/SB0/n25 ), .B0(\U1/aes_core/SB0/n21 ), .Y(
        \U1/aes_core/SB0/n1380 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1146  ( .A(\U1/aes_core/SB0/n1345 ), .B(
        \U1/aes_core/SB0/n52 ), .Y(\U1/aes_core/SB0/n13 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1145  ( .A0(\U1/aes_core/SB0/n47 ), .A1(
        \U1/aes_core/SB0/n13 ), .B0(\U1/aes_core/SB0/n1308 ), .B1(
        \U1/aes_core/SB0/n49 ), .Y(\U1/aes_core/SB0/n1381 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U1144  ( .A0(\U1/aes_core/SB0/n1379 ), 
        .A1(\U1/aes_core/SB0/n1323 ), .B0(\U1/aes_core/SB0/n1380 ), .C0(
        \U1/aes_core/SB0/n1381 ), .Y(\U1/aes_core/SB0/n1378 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1143  ( .A(\U1/aes_core/SB0/n1361 ), .B(
        \U1/aes_core/SB0/n1374 ), .C(\U1/aes_core/SB0/n1375 ), .D(
        \U1/aes_core/SB0/n1376 ), .E(\U1/aes_core/SB0/n1377 ), .F(
        \U1/aes_core/SB0/n1378 ), .Y(\U1/aes_core/sb0 [13]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1142  ( .A0(\U1/aes_core/SB0/n11 ), 
        .A1(\U1/aes_core/SB0/n58 ), .B0(\U1/aes_core/SB0/n53 ), .B1(
        \U1/aes_core/SB0/n1292 ), .C0(\U1/aes_core/SB0/n1373 ), .Y(
        \U1/aes_core/SB0/n1364 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1141  ( .A0(\U1/aes_core/SB0/n79 ), .A1(
        \U1/aes_core/SB0/n1294 ), .B0(\U1/aes_core/SB0/n32 ), .Y(
        \U1/aes_core/SB0/n1369 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1140  ( .A0(\U1/aes_core/SB0/n1307 ), 
        .A1(\U1/aes_core/SB0/n55 ), .B0(\U1/aes_core/SB0/n1302 ), .Y(
        \U1/aes_core/SB0/n1370 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1139  ( .A(\U1/aes_core/SB0/n1352 ), .B(
        \U1/aes_core/SB0/n8 ), .Y(\U1/aes_core/SB0/n26 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1138  ( .A0(\U1/aes_core/SB0/n49 ), .A1(
        \U1/aes_core/SB0/n86 ), .B0(\U1/aes_core/SB0/n26 ), .Y(
        \U1/aes_core/SB0/n1371 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1137  ( .A(\U1/aes_core/SB0/n1369 ), .B(
        \U1/aes_core/SB0/n1370 ), .C(\U1/aes_core/SB0/n1371 ), .D(
        \U1/aes_core/SB0/n1372 ), .Y(\U1/aes_core/SB0/n1365 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1136  ( .A(\U1/aes_core/SB0/n11 ), .B(
        \U1/aes_core/SB0/n10 ), .Y(\U1/aes_core/SB0/n1296 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1135  ( .A(\U1/aes_core/SB0/n22 ), .B(
        \U1/aes_core/SB0/n1296 ), .Y(\U1/aes_core/SB0/n1368 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1134  ( .A0(\U1/aes_core/SB0/n1305 ), 
        .A1(\U1/aes_core/SB0/n1367 ), .B0(\U1/aes_core/SB0/n1368 ), .B1(
        \U1/aes_core/SB0/n1352 ), .C0(\U1/aes_core/SB0/n1354 ), .C1(
        \U1/aes_core/SB0/n1323 ), .Y(\U1/aes_core/SB0/n1366 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1133  ( .A(\U1/aes_core/SB0/n1361 ), .B(
        \U1/aes_core/SB0/n1362 ), .C(\U1/aes_core/SB0/n1363 ), .D(
        \U1/aes_core/SB0/n1364 ), .E(\U1/aes_core/SB0/n1365 ), .F(
        \U1/aes_core/SB0/n1366 ), .Y(\U1/aes_core/sb0 [14]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1132  ( .A0(\U1/aes_core/SB0/n1360 ), 
        .A1(\U1/aes_core/SB0/n52 ), .B0(\U1/aes_core/SB0/n1292 ), .Y(
        \U1/aes_core/SB0/n1348 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U1131  ( .A(\U1/aes_core/SB0/n1357 ), .B(
        \U1/aes_core/SB0/n1358 ), .C(\U1/aes_core/SB0/n1359 ), .Y(
        \U1/aes_core/SB0/n1349 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U1130  ( .A(\U1/aes_core/SB0/n1308 ), .B(
        \U1/aes_core/SB0/n1304 ), .C(\U1/aes_core/SB0/n72 ), .Y(
        \U1/aes_core/SB0/n1355 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1129  ( .A0(\U1/aes_core/SB0/n1353 ), 
        .A1(\U1/aes_core/SB0/n1354 ), .B0(\U1/aes_core/SB0/n1355 ), .B1(
        \U1/aes_core/SB0/n1297 ), .C0(\U1/aes_core/SB0/n1356 ), .C1(
        \U1/aes_core/SB0/n74 ), .Y(\U1/aes_core/SB0/n1350 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U1128  ( .A0(\U1/aes_core/SB0/n11 ), .A1(
        \U1/aes_core/SB0/n1323 ), .B0(\U1/aes_core/SB0/n10 ), .B1(
        \U1/aes_core/SB0/n1352 ), .Y(\U1/aes_core/SB0/n1351 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1127  ( .A(\U1/aes_core/SB0/n1346 ), .B(
        \U1/aes_core/SB0/n1347 ), .C(\U1/aes_core/SB0/n1348 ), .D(
        \U1/aes_core/SB0/n1349 ), .E(\U1/aes_core/SB0/n1350 ), .F(
        \U1/aes_core/SB0/n1351 ), .Y(\U1/aes_core/SB0/n2 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U1126  ( .A0(\U1/aes_core/SB0/n76 ), .A1(
        \U1/aes_core/SB0/n7 ), .B0(\U1/aes_core/SB0/n1345 ), .Y(
        \U1/aes_core/SB0/n1329 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB0/U1125  ( .A0(\U1/aes_core/SB0/n1343 ), 
        .A1(\U1/aes_core/SB0/n85 ), .B0(\U1/aes_core/SB0/n1344 ), .B1(
        \U1/aes_core/SB0/n25 ), .Y(\U1/aes_core/SB0/n1330 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1124  ( .A0(\U1/aes_core/SB0/n73 ), 
        .A1(\U1/aes_core/SB0/n10 ), .B0(\U1/aes_core/SB0/n1341 ), .B1(
        \U1/aes_core/SB0/n1342 ), .C0(\U1/aes_core/SB0/n1323 ), .C1(
        \U1/aes_core/SB0/n1297 ), .Y(\U1/aes_core/SB0/n1331 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1123  ( .A(\U1/aes_core/SB0/n1337 ), .B(
        \U1/aes_core/SB0/n1338 ), .C(\U1/aes_core/SB0/n1339 ), .D(
        \U1/aes_core/SB0/n1340 ), .Y(\U1/aes_core/SB0/n1332 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1122  ( .AN(\U1/aes_core/SB0/n1334 ), 
        .B(\U1/aes_core/SB0/n1335 ), .C(\U1/aes_core/SB0/n1336 ), .Y(
        \U1/aes_core/SB0/n1333 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1121  ( .A(\U1/aes_core/SB0/n1328 ), .B(
        \U1/aes_core/SB0/n1329 ), .C(\U1/aes_core/SB0/n1330 ), .D(
        \U1/aes_core/SB0/n1331 ), .E(\U1/aes_core/SB0/n1332 ), .F(
        \U1/aes_core/SB0/n1333 ), .Y(\U1/aes_core/SB0/n60 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1120  ( .A0(\U1/aes_core/SB0/n47 ), .A1(
        \U1/aes_core/SB0/n27 ), .B0(\U1/aes_core/SB0/n1308 ), .Y(
        \U1/aes_core/SB0/n1324 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1119  ( .A(\U1/aes_core/SB0/n1324 ), .B(
        \U1/aes_core/SB0/n1325 ), .C(\U1/aes_core/SB0/n1326 ), .D(
        \U1/aes_core/SB0/n1327 ), .Y(\U1/aes_core/SB0/n1311 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1118  ( .A0(\U1/aes_core/SB0/n53 ), 
        .A1(\U1/aes_core/SB0/n1292 ), .B0(\U1/aes_core/SB0/n75 ), .B1(
        \U1/aes_core/SB0/n74 ), .C0(\U1/aes_core/SB0/n45 ), .C1(
        \U1/aes_core/SB0/n1323 ), .Y(\U1/aes_core/SB0/n1312 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1117  ( .A(\U1/aes_core/SB0/n1319 ), .B(
        \U1/aes_core/SB0/n1320 ), .C(\U1/aes_core/SB0/n1321 ), .D(
        \U1/aes_core/SB0/n1322 ), .Y(\U1/aes_core/SB0/n1313 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U1116  ( .A(\U1/aes_core/SB0/n1315 ), .B(
        \U1/aes_core/SB0/n1316 ), .C(\U1/aes_core/SB0/n1317 ), .D(
        \U1/aes_core/SB0/n1318 ), .Y(\U1/aes_core/SB0/n1314 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1115  ( .A(\U1/aes_core/SB0/n1311 ), .B(
        \U1/aes_core/SB0/n1312 ), .C(\U1/aes_core/SB0/n1313 ), .D(
        \U1/aes_core/SB0/n1314 ), .Y(\U1/aes_core/SB0/n1310 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1114  ( .A(\U1/aes_core/SB0/n1310 ), .Y(
        \U1/aes_core/SB0/n69 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1113  ( .A0(\U1/aes_core/SB0/n1307 ), 
        .A1(\U1/aes_core/SB0/n24 ), .B0(\U1/aes_core/SB0/n1308 ), .B1(
        \U1/aes_core/SB0/n1309 ), .Y(\U1/aes_core/SB0/n1306 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U1112  ( .A0(\U1/aes_core/SB0/n1305 ), 
        .A1(\U1/aes_core/SB0/n45 ), .B0(\U1/aes_core/SB0/n69 ), .C0(
        \U1/aes_core/SB0/n1306 ), .Y(\U1/aes_core/SB0/n1289 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U1111  ( .A1N(\U1/aes_core/SB0/n1303 ), 
        .A0(\U1/aes_core/SB0/n1304 ), .B0(\U1/aes_core/SB0/n22 ), .Y(
        \U1/aes_core/SB0/n1299 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1110  ( .A0(\U1/aes_core/SB0/n27 ), .A1(
        \U1/aes_core/SB0/n32 ), .B0(\U1/aes_core/SB0/n1302 ), .Y(
        \U1/aes_core/SB0/n1300 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1109  ( .AN(\U1/aes_core/SB0/n1298 ), 
        .B(\U1/aes_core/SB0/n1299 ), .C(\U1/aes_core/SB0/n1300 ), .D(
        \U1/aes_core/SB0/n1301 ), .Y(\U1/aes_core/SB0/n1290 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1108  ( .A(\U1/aes_core/SB0/n1297 ), .B(
        \U1/aes_core/SB0/n11 ), .Y(\U1/aes_core/SB0/n1295 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1107  ( .A0(\U1/aes_core/SB0/n1294 ), 
        .A1(\U1/aes_core/SB0/n1295 ), .B0(\U1/aes_core/SB0/n72 ), .B1(
        \U1/aes_core/SB0/n1296 ), .Y(\U1/aes_core/SB0/n1293 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1106  ( .A0(\U1/aes_core/SB0/n73 ), 
        .A1(\U1/aes_core/SB0/n7 ), .B0(\U1/aes_core/SB0/n1292 ), .B1(
        \U1/aes_core/SB0/n12 ), .C0(\U1/aes_core/SB0/n1293 ), .Y(
        \U1/aes_core/SB0/n1291 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U1105  ( .A(\U1/aes_core/SB0/n2 ), .B(
        \U1/aes_core/SB0/n60 ), .C(\U1/aes_core/SB0/n1288 ), .D(
        \U1/aes_core/SB0/n1289 ), .E(\U1/aes_core/SB0/n1290 ), .F(
        \U1/aes_core/SB0/n1291 ), .Y(\U1/aes_core/sb0 [15]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1104  ( .A(Dout[119]), .B(Dout[118]), .Y(
        \U1/aes_core/SB0/n1269 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1103  ( .A(Dout[117]), .B(Dout[116]), .Y(
        \U1/aes_core/SB0/n1278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1102  ( .A(\U1/aes_core/SB0/n1269 ), .B(
        \U1/aes_core/SB0/n1278 ), .Y(\U1/aes_core/SB0/n1204 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1101  ( .A(Dout[113]), .Y(
        \U1/aes_core/SB0/n1284 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1100  ( .A(Dout[112]), .Y(
        \U1/aes_core/SB0/n1287 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1099  ( .A(\U1/aes_core/SB0/n1284 ), .B(
        \U1/aes_core/SB0/n1287 ), .Y(\U1/aes_core/SB0/n1277 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1098  ( .A(Dout[115]), .B(Dout[114]), .Y(
        \U1/aes_core/SB0/n1257 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1097  ( .A(\U1/aes_core/SB0/n1277 ), .B(
        \U1/aes_core/SB0/n1257 ), .Y(\U1/aes_core/SB0/n894 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1096  ( .A(\U1/aes_core/SB0/n1204 ), .B(
        \U1/aes_core/SB0/n894 ), .Y(\U1/aes_core/SB0/n1113 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U1095  ( .A(Dout[114]), .B(Dout[115]), .Y(
        \U1/aes_core/SB0/n1274 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1094  ( .A(\U1/aes_core/SB0/n1274 ), .B(
        \U1/aes_core/SB0/n1277 ), .Y(\U1/aes_core/SB0/n956 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1093  ( .A(Dout[119]), .Y(
        \U1/aes_core/SB0/n1281 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1092  ( .A(\U1/aes_core/SB0/n1281 ), .B(
        Dout[118]), .Y(\U1/aes_core/SB0/n1251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1091  ( .A(\U1/aes_core/SB0/n1251 ), .B(
        \U1/aes_core/SB0/n1278 ), .Y(\U1/aes_core/SB0/n1205 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1090  ( .A(\U1/aes_core/SB0/n956 ), .B(
        \U1/aes_core/SB0/n1205 ), .Y(\U1/aes_core/SB0/n990 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1089  ( .A(Dout[115]), .Y(
        \U1/aes_core/SB0/n1286 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U1088  ( .A(Dout[114]), .B(
        \U1/aes_core/SB0/n1286 ), .Y(\U1/aes_core/SB0/n1276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1087  ( .A(\U1/aes_core/SB0/n1277 ), .B(
        \U1/aes_core/SB0/n1276 ), .Y(\U1/aes_core/SB0/n1051 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1086  ( .A(\U1/aes_core/SB0/n1051 ), .Y(
        \U1/aes_core/SB0/n860 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1085  ( .A(Dout[116]), .Y(
        \U1/aes_core/SB0/n1285 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1084  ( .A(\U1/aes_core/SB0/n1285 ), .B(
        Dout[117]), .Y(\U1/aes_core/SB0/n1270 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1083  ( .A(Dout[118]), .Y(
        \U1/aes_core/SB0/n1282 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1082  ( .A(\U1/aes_core/SB0/n1282 ), .B(
        Dout[119]), .Y(\U1/aes_core/SB0/n1260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1081  ( .A(\U1/aes_core/SB0/n1270 ), .B(
        \U1/aes_core/SB0/n1260 ), .Y(\U1/aes_core/SB0/n1004 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1080  ( .A(\U1/aes_core/SB0/n1004 ), .Y(
        \U1/aes_core/SB0/n906 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1079  ( .A(\U1/aes_core/SB0/n860 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1073 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1078  ( .A(\U1/aes_core/SB0/n1204 ), .Y(
        \U1/aes_core/SB0/n891 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1077  ( .A(Dout[113]), .B(Dout[112]), .Y(
        \U1/aes_core/SB0/n1273 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1076  ( .A(\U1/aes_core/SB0/n1273 ), .B(
        \U1/aes_core/SB0/n1257 ), .Y(\U1/aes_core/SB0/n938 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1075  ( .A(\U1/aes_core/SB0/n938 ), .Y(
        \U1/aes_core/SB0/n850 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1074  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n850 ), .Y(\U1/aes_core/SB0/n933 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1073  ( .A(\U1/aes_core/SB0/n1287 ), .B(
        Dout[113]), .Y(\U1/aes_core/SB0/n1258 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1072  ( .A(\U1/aes_core/SB0/n1276 ), .B(
        \U1/aes_core/SB0/n1258 ), .Y(\U1/aes_core/SB0/n1064 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1071  ( .A(\U1/aes_core/SB0/n1064 ), .Y(
        \U1/aes_core/SB0/n949 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1070  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1095 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U1069  ( .A(\U1/aes_core/SB0/n1073 ), .B(
        \U1/aes_core/SB0/n933 ), .C(\U1/aes_core/SB0/n1095 ), .Y(
        \U1/aes_core/SB0/n1238 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1068  ( .A(\U1/aes_core/SB0/n1278 ), .B(
        \U1/aes_core/SB0/n1260 ), .Y(\U1/aes_core/SB0/n1005 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1067  ( .A(\U1/aes_core/SB0/n1286 ), .B(
        Dout[114]), .Y(\U1/aes_core/SB0/n1267 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1066  ( .A(\U1/aes_core/SB0/n1267 ), .B(
        \U1/aes_core/SB0/n1258 ), .Y(\U1/aes_core/SB0/n1007 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1065  ( .A(\U1/aes_core/SB0/n1005 ), .B(
        \U1/aes_core/SB0/n1007 ), .Y(\U1/aes_core/SB0/n1118 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1064  ( .A(\U1/aes_core/SB0/n1205 ), .Y(
        \U1/aes_core/SB0/n889 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1063  ( .A(Dout[117]), .Y(
        \U1/aes_core/SB0/n1283 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1062  ( .A(\U1/aes_core/SB0/n1285 ), .B(
        \U1/aes_core/SB0/n1283 ), .Y(\U1/aes_core/SB0/n1259 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1061  ( .A(\U1/aes_core/SB0/n1269 ), .B(
        \U1/aes_core/SB0/n1259 ), .Y(\U1/aes_core/SB0/n846 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1060  ( .A(\U1/aes_core/SB0/n846 ), .Y(
        \U1/aes_core/SB0/n915 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1059  ( .A(\U1/aes_core/SB0/n1284 ), .B(
        Dout[112]), .Y(\U1/aes_core/SB0/n1268 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1058  ( .A(\U1/aes_core/SB0/n1268 ), .B(
        \U1/aes_core/SB0/n1257 ), .Y(\U1/aes_core/SB0/n881 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1057  ( .A(\U1/aes_core/SB0/n881 ), .Y(
        \U1/aes_core/SB0/n1059 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1056  ( .A0(\U1/aes_core/SB0/n889 ), 
        .A1(\U1/aes_core/SB0/n915 ), .B0(\U1/aes_core/SB0/n1059 ), .Y(
        \U1/aes_core/SB0/n1279 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1055  ( .A(\U1/aes_core/SB0/n1273 ), .B(
        \U1/aes_core/SB0/n1276 ), .Y(\U1/aes_core/SB0/n893 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1054  ( .A(\U1/aes_core/SB0/n893 ), .Y(
        \U1/aes_core/SB0/n907 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1053  ( .A(\U1/aes_core/SB0/n1283 ), .B(
        Dout[116]), .Y(\U1/aes_core/SB0/n1252 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1052  ( .A(\U1/aes_core/SB0/n1260 ), .B(
        \U1/aes_core/SB0/n1252 ), .Y(\U1/aes_core/SB0/n853 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1051  ( .A(\U1/aes_core/SB0/n1005 ), .B(
        \U1/aes_core/SB0/n853 ), .Y(\U1/aes_core/SB0/n1140 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1050  ( .A(\U1/aes_core/SB0/n1281 ), .B(
        \U1/aes_core/SB0/n1282 ), .Y(\U1/aes_core/SB0/n1261 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1049  ( .A(\U1/aes_core/SB0/n1270 ), .B(
        \U1/aes_core/SB0/n1261 ), .Y(\U1/aes_core/SB0/n878 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1048  ( .A(\U1/aes_core/SB0/n878 ), .Y(
        \U1/aes_core/SB0/n1160 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1047  ( .A0(\U1/aes_core/SB0/n907 ), 
        .A1(\U1/aes_core/SB0/n1140 ), .B0(\U1/aes_core/SB0/n1160 ), .B1(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1280 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U1046  ( .AN(\U1/aes_core/SB0/n1118 ), 
        .B(\U1/aes_core/SB0/n1279 ), .C(\U1/aes_core/SB0/n1280 ), .Y(
        \U1/aes_core/SB0/n1239 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1045  ( .A(\U1/aes_core/SB0/n1278 ), .B(
        \U1/aes_core/SB0/n1261 ), .Y(\U1/aes_core/SB0/n988 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1044  ( .A(\U1/aes_core/SB0/n1274 ), .B(
        \U1/aes_core/SB0/n1273 ), .Y(\U1/aes_core/SB0/n843 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1043  ( .A(\U1/aes_core/SB0/n1251 ), .B(
        \U1/aes_core/SB0/n1270 ), .Y(\U1/aes_core/SB0/n937 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1042  ( .A(\U1/aes_core/SB0/n1274 ), .B(
        \U1/aes_core/SB0/n1268 ), .Y(\U1/aes_core/SB0/n940 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1041  ( .A(\U1/aes_core/SB0/n1277 ), .B(
        \U1/aes_core/SB0/n1267 ), .Y(\U1/aes_core/SB0/n935 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1040  ( .A(\U1/aes_core/SB0/n935 ), .Y(
        \U1/aes_core/SB0/n955 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1039  ( .A(\U1/aes_core/SB0/n853 ), .Y(
        \U1/aes_core/SB0/n1145 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1038  ( .A(\U1/aes_core/SB0/n1276 ), .B(
        \U1/aes_core/SB0/n1268 ), .Y(\U1/aes_core/SB0/n917 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1037  ( .A(\U1/aes_core/SB0/n917 ), .Y(
        \U1/aes_core/SB0/n892 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U1036  ( .A0(\U1/aes_core/SB0/n955 ), 
        .A1(\U1/aes_core/SB0/n891 ), .B0(\U1/aes_core/SB0/n1145 ), .B1(
        \U1/aes_core/SB0/n892 ), .Y(\U1/aes_core/SB0/n1275 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U1035  ( .A0(\U1/aes_core/SB0/n988 ), 
        .A1(\U1/aes_core/SB0/n843 ), .B0(\U1/aes_core/SB0/n937 ), .B1(
        \U1/aes_core/SB0/n940 ), .C0(\U1/aes_core/SB0/n1275 ), .Y(
        \U1/aes_core/SB0/n1240 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1034  ( .A(\U1/aes_core/SB0/n935 ), .B(
        \U1/aes_core/SB0/n988 ), .Y(\U1/aes_core/SB0/n1152 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1033  ( .A(\U1/aes_core/SB0/n940 ), .B(
        \U1/aes_core/SB0/n1005 ), .Y(\U1/aes_core/SB0/n1142 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1032  ( .A(\U1/aes_core/SB0/n1142 ), .Y(
        \U1/aes_core/SB0/n1271 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1031  ( .A(\U1/aes_core/SB0/n1274 ), .B(
        \U1/aes_core/SB0/n1258 ), .Y(\U1/aes_core/SB0/n865 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1030  ( .A(\U1/aes_core/SB0/n865 ), .Y(
        \U1/aes_core/SB0/n916 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1029  ( .A(\U1/aes_core/SB0/n1273 ), .B(
        \U1/aes_core/SB0/n1267 ), .Y(\U1/aes_core/SB0/n880 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1028  ( .A(\U1/aes_core/SB0/n880 ), .Y(
        \U1/aes_core/SB0/n869 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U1027  ( .A0(\U1/aes_core/SB0/n916 ), 
        .A1(\U1/aes_core/SB0/n869 ), .B0(\U1/aes_core/SB0/n915 ), .Y(
        \U1/aes_core/SB0/n1272 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1026  ( .A(\U1/aes_core/SB0/n1269 ), .B(
        \U1/aes_core/SB0/n1252 ), .Y(\U1/aes_core/SB0/n864 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1025  ( .A(\U1/aes_core/SB0/n864 ), .Y(
        \U1/aes_core/SB0/n914 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1024  ( .A(\U1/aes_core/SB0/n914 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1125 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1023  ( .AN(\U1/aes_core/SB0/n1152 ), 
        .B(\U1/aes_core/SB0/n1271 ), .C(\U1/aes_core/SB0/n1272 ), .D(
        \U1/aes_core/SB0/n1125 ), .Y(\U1/aes_core/SB0/n1262 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1022  ( .A(\U1/aes_core/SB0/n1259 ), .B(
        \U1/aes_core/SB0/n1261 ), .Y(\U1/aes_core/SB0/n844 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1021  ( .A(\U1/aes_core/SB0/n1269 ), .B(
        \U1/aes_core/SB0/n1270 ), .Y(\U1/aes_core/SB0/n852 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U1020  ( .A0(\U1/aes_core/SB0/n1205 ), 
        .A1(\U1/aes_core/SB0/n1051 ), .B0(\U1/aes_core/SB0/n844 ), .B1(
        \U1/aes_core/SB0/n935 ), .C0(\U1/aes_core/SB0/n852 ), .C1(
        \U1/aes_core/SB0/n917 ), .Y(\U1/aes_core/SB0/n1263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1019  ( .A(\U1/aes_core/SB0/n893 ), .B(
        \U1/aes_core/SB0/n1205 ), .Y(\U1/aes_core/SB0/n1067 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1018  ( .A(\U1/aes_core/SB0/n1145 ), .B(
        \U1/aes_core/SB0/n955 ), .Y(\U1/aes_core/SB0/n1114 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1017  ( .A(\U1/aes_core/SB0/n892 ), .B(
        \U1/aes_core/SB0/n891 ), .Y(\U1/aes_core/SB0/n1094 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1016  ( .A(\U1/aes_core/SB0/n937 ), .Y(
        \U1/aes_core/SB0/n863 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1015  ( .A(\U1/aes_core/SB0/n863 ), .B(
        \U1/aes_core/SB0/n1059 ), .Y(\U1/aes_core/SB0/n1056 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1014  ( .AN(\U1/aes_core/SB0/n1067 ), 
        .B(\U1/aes_core/SB0/n1114 ), .C(\U1/aes_core/SB0/n1094 ), .D(
        \U1/aes_core/SB0/n1056 ), .Y(\U1/aes_core/SB0/n1264 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1013  ( .A(\U1/aes_core/SB0/n1251 ), .B(
        \U1/aes_core/SB0/n1259 ), .Y(\U1/aes_core/SB0/n1144 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1012  ( .A(\U1/aes_core/SB0/n1144 ), .B(
        \U1/aes_core/SB0/n881 ), .Y(\U1/aes_core/SB0/n964 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1011  ( .A(\U1/aes_core/SB0/n1267 ), .B(
        \U1/aes_core/SB0/n1268 ), .Y(\U1/aes_core/SB0/n845 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1010  ( .A(\U1/aes_core/SB0/n878 ), .B(
        \U1/aes_core/SB0/n845 ), .Y(\U1/aes_core/SB0/n999 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1009  ( .A(\U1/aes_core/SB0/n999 ), .Y(
        \U1/aes_core/SB0/n1266 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1008  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n1059 ), .Y(\U1/aes_core/SB0/n980 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1007  ( .A(\U1/aes_core/SB0/n845 ), .Y(
        \U1/aes_core/SB0/n862 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1006  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n862 ), .Y(\U1/aes_core/SB0/n929 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U1005  ( .AN(\U1/aes_core/SB0/n964 ), 
        .B(\U1/aes_core/SB0/n1266 ), .C(\U1/aes_core/SB0/n980 ), .D(
        \U1/aes_core/SB0/n929 ), .Y(\U1/aes_core/SB0/n1265 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U1004  ( .A(\U1/aes_core/SB0/n1262 ), .B(
        \U1/aes_core/SB0/n1263 ), .C(\U1/aes_core/SB0/n1264 ), .D(
        \U1/aes_core/SB0/n1265 ), .Y(\U1/aes_core/SB0/n1164 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1003  ( .A(\U1/aes_core/SB0/n938 ), .B(
        \U1/aes_core/SB0/n1144 ), .Y(\U1/aes_core/SB0/n930 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U1002  ( .A(\U1/aes_core/SB0/n1252 ), .B(
        \U1/aes_core/SB0/n1261 ), .Y(\U1/aes_core/SB0/n1048 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U1001  ( .A(\U1/aes_core/SB0/n956 ), .B(
        \U1/aes_core/SB0/n1048 ), .Y(\U1/aes_core/SB0/n1077 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U1000  ( .A(\U1/aes_core/SB0/n844 ), .Y(
        \U1/aes_core/SB0/n888 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U999  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n907 ), .Y(\U1/aes_core/SB0/n1128 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U998  ( .A0(\U1/aes_core/SB0/n1048 ), 
        .A1(\U1/aes_core/SB0/n845 ), .B0(\U1/aes_core/SB0/n1128 ), .Y(
        \U1/aes_core/SB0/n1253 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U997  ( .A(\U1/aes_core/SB0/n1007 ), .Y(
        \U1/aes_core/SB0/n912 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U996  ( .A(\U1/aes_core/SB0/n912 ), .B(
        \U1/aes_core/SB0/n889 ), .Y(\U1/aes_core/SB0/n911 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U995  ( .A(\U1/aes_core/SB0/n889 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n952 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U994  ( .A(\U1/aes_core/SB0/n1259 ), .B(
        \U1/aes_core/SB0/n1260 ), .Y(\U1/aes_core/SB0/n882 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U993  ( .A(\U1/aes_core/SB0/n882 ), .Y(
        \U1/aes_core/SB0/n1133 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U992  ( .A(\U1/aes_core/SB0/n916 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n1109 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U991  ( .A(\U1/aes_core/SB0/n894 ), .Y(
        \U1/aes_core/SB0/n913 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U990  ( .A(\U1/aes_core/SB0/n913 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n1045 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U989  ( .A(\U1/aes_core/SB0/n911 ), .B(
        \U1/aes_core/SB0/n952 ), .C(\U1/aes_core/SB0/n1109 ), .D(
        \U1/aes_core/SB0/n1045 ), .Y(\U1/aes_core/SB0/n1254 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U988  ( .A(\U1/aes_core/SB0/n892 ), .B(
        \U1/aes_core/SB0/n914 ), .Y(\U1/aes_core/SB0/n985 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U987  ( .A(\U1/aes_core/SB0/n850 ), .B(
        \U1/aes_core/SB0/n914 ), .Y(\U1/aes_core/SB0/n994 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U986  ( .A(\U1/aes_core/SB0/n852 ), .Y(
        \U1/aes_core/SB0/n859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U985  ( .A(\U1/aes_core/SB0/n955 ), .B(
        \U1/aes_core/SB0/n859 ), .Y(\U1/aes_core/SB0/n1148 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U984  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n916 ), .Y(\U1/aes_core/SB0/n1011 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U983  ( .A(\U1/aes_core/SB0/n985 ), .B(
        \U1/aes_core/SB0/n994 ), .C(\U1/aes_core/SB0/n1148 ), .D(
        \U1/aes_core/SB0/n1011 ), .Y(\U1/aes_core/SB0/n1255 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U982  ( .A(\U1/aes_core/SB0/n940 ), .Y(
        \U1/aes_core/SB0/n971 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U981  ( .A(\U1/aes_core/SB0/n1145 ), .B(
        \U1/aes_core/SB0/n971 ), .Y(\U1/aes_core/SB0/n1162 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U980  ( .A(\U1/aes_core/SB0/n1257 ), .B(
        \U1/aes_core/SB0/n1258 ), .Y(\U1/aes_core/SB0/n905 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U979  ( .A(\U1/aes_core/SB0/n905 ), .Y(
        \U1/aes_core/SB0/n871 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U978  ( .A(\U1/aes_core/SB0/n1145 ), .B(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n1097 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U977  ( .A(\U1/aes_core/SB0/n956 ), .Y(
        \U1/aes_core/SB0/n848 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U976  ( .A(\U1/aes_core/SB0/n848 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1062 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U975  ( .A(\U1/aes_core/SB0/n915 ), .B(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n887 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U974  ( .A(\U1/aes_core/SB0/n1162 ), .B(
        \U1/aes_core/SB0/n1097 ), .C(\U1/aes_core/SB0/n1062 ), .D(
        \U1/aes_core/SB0/n887 ), .Y(\U1/aes_core/SB0/n1256 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U973  ( .A(\U1/aes_core/SB0/n930 ), .B(
        \U1/aes_core/SB0/n1077 ), .C(\U1/aes_core/SB0/n1253 ), .D(
        \U1/aes_core/SB0/n1254 ), .E(\U1/aes_core/SB0/n1255 ), .F(
        \U1/aes_core/SB0/n1256 ), .Y(\U1/aes_core/SB0/n1175 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U972  ( .A(\U1/aes_core/SB0/n1175 ), .Y(
        \U1/aes_core/SB0/n1242 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U971  ( .A(\U1/aes_core/SB0/n880 ), .B(
        \U1/aes_core/SB0/n1048 ), .Y(\U1/aes_core/SB0/n1151 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U970  ( .A(\U1/aes_core/SB0/n1251 ), .B(
        \U1/aes_core/SB0/n1252 ), .Y(\U1/aes_core/SB0/n883 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U969  ( .A(\U1/aes_core/SB0/n883 ), .B(
        \U1/aes_core/SB0/n1007 ), .Y(\U1/aes_core/SB0/n998 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U968  ( .A(\U1/aes_core/SB0/n998 ), .Y(
        \U1/aes_core/SB0/n1249 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U967  ( .A(\U1/aes_core/SB0/n1005 ), .Y(
        \U1/aes_core/SB0/n858 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U966  ( .A0(\U1/aes_core/SB0/n1133 ), 
        .A1(\U1/aes_core/SB0/n858 ), .B0(\U1/aes_core/SB0/n871 ), .Y(
        \U1/aes_core/SB0/n1250 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U965  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n971 ), .Y(\U1/aes_core/SB0/n1126 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U964  ( .AN(\U1/aes_core/SB0/n1151 ), 
        .B(\U1/aes_core/SB0/n1249 ), .C(\U1/aes_core/SB0/n1250 ), .D(
        \U1/aes_core/SB0/n1126 ), .Y(\U1/aes_core/SB0/n1245 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U963  ( .A0(\U1/aes_core/SB0/n894 ), 
        .A1(\U1/aes_core/SB0/n846 ), .B0(\U1/aes_core/SB0/n988 ), .B1(
        \U1/aes_core/SB0/n940 ), .C0(\U1/aes_core/SB0/n881 ), .C1(
        \U1/aes_core/SB0/n864 ), .Y(\U1/aes_core/SB0/n1246 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U962  ( .A(\U1/aes_core/SB0/n846 ), .B(
        \U1/aes_core/SB0/n843 ), .Y(\U1/aes_core/SB0/n1086 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U961  ( .A(\U1/aes_core/SB0/n858 ), .B(
        \U1/aes_core/SB0/n916 ), .Y(\U1/aes_core/SB0/n927 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U960  ( .A(\U1/aes_core/SB0/n955 ), .B(
        \U1/aes_core/SB0/n858 ), .Y(\U1/aes_core/SB0/n993 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U959  ( .A(\U1/aes_core/SB0/n971 ), .B(
        \U1/aes_core/SB0/n891 ), .Y(\U1/aes_core/SB0/n1147 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U958  ( .AN(\U1/aes_core/SB0/n1086 ), 
        .B(\U1/aes_core/SB0/n927 ), .C(\U1/aes_core/SB0/n993 ), .D(
        \U1/aes_core/SB0/n1147 ), .Y(\U1/aes_core/SB0/n1247 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U957  ( .A(\U1/aes_core/SB0/n848 ), .B(
        \U1/aes_core/SB0/n863 ), .Y(\U1/aes_core/SB0/n1074 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U956  ( .A(\U1/aes_core/SB0/n971 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n981 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U955  ( .A(\U1/aes_core/SB0/n1145 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1106 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U954  ( .A(\U1/aes_core/SB0/n912 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1061 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U953  ( .A(\U1/aes_core/SB0/n1074 ), .B(
        \U1/aes_core/SB0/n981 ), .C(\U1/aes_core/SB0/n1106 ), .D(
        \U1/aes_core/SB0/n1061 ), .Y(\U1/aes_core/SB0/n1248 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U952  ( .A(\U1/aes_core/SB0/n1245 ), .B(
        \U1/aes_core/SB0/n1246 ), .C(\U1/aes_core/SB0/n1247 ), .D(
        \U1/aes_core/SB0/n1248 ), .Y(\U1/aes_core/SB0/n1244 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U951  ( .A(\U1/aes_core/SB0/n1244 ), .Y(
        \U1/aes_core/SB0/n866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U950  ( .A(\U1/aes_core/SB0/n850 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1243 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U949  ( .AN(\U1/aes_core/SB0/n1164 ), 
        .B(\U1/aes_core/SB0/n1242 ), .C(\U1/aes_core/SB0/n866 ), .D(
        \U1/aes_core/SB0/n1243 ), .Y(\U1/aes_core/SB0/n1241 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U948  ( .A(\U1/aes_core/SB0/n1113 ), .B(
        \U1/aes_core/SB0/n990 ), .C(\U1/aes_core/SB0/n1238 ), .D(
        \U1/aes_core/SB0/n1239 ), .E(\U1/aes_core/SB0/n1240 ), .F(
        \U1/aes_core/SB0/n1241 ), .Y(\U1/aes_core/SB0/n1185 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U947  ( .A(\U1/aes_core/SB0/n865 ), .B(
        \U1/aes_core/SB0/n1205 ), .Y(\U1/aes_core/SB0/n1068 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U946  ( .A(\U1/aes_core/SB0/n915 ), .B(
        \U1/aes_core/SB0/n848 ), .Y(\U1/aes_core/SB0/n991 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U945  ( .A(\U1/aes_core/SB0/n859 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1115 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U944  ( .A(\U1/aes_core/SB0/n1144 ), .Y(
        \U1/aes_core/SB0/n870 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U943  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1092 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U942  ( .AN(\U1/aes_core/SB0/n1068 ), 
        .B(\U1/aes_core/SB0/n991 ), .C(\U1/aes_core/SB0/n1115 ), .D(
        \U1/aes_core/SB0/n1092 ), .Y(\U1/aes_core/SB0/n1231 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U941  ( .A(\U1/aes_core/SB0/n878 ), .B(
        \U1/aes_core/SB0/n1007 ), .Y(\U1/aes_core/SB0/n965 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U940  ( .A(\U1/aes_core/SB0/n955 ), .B(
        \U1/aes_core/SB0/n889 ), .Y(\U1/aes_core/SB0/n1135 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U939  ( .A0(\U1/aes_core/SB0/n869 ), .A1(
        \U1/aes_core/SB0/n949 ), .B0(\U1/aes_core/SB0/n1145 ), .Y(
        \U1/aes_core/SB0/n1237 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U938  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1043 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U937  ( .AN(\U1/aes_core/SB0/n965 ), .B(
        \U1/aes_core/SB0/n1135 ), .C(\U1/aes_core/SB0/n1237 ), .D(
        \U1/aes_core/SB0/n1043 ), .Y(\U1/aes_core/SB0/n1236 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U936  ( .A(\U1/aes_core/SB0/n1236 ), .Y(
        \U1/aes_core/SB0/n1232 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U935  ( .A(\U1/aes_core/SB0/n988 ), .Y(
        \U1/aes_core/SB0/n868 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U934  ( .A(\U1/aes_core/SB0/n843 ), .Y(
        \U1/aes_core/SB0/n948 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U933  ( .A0(\U1/aes_core/SB0/n848 ), 
        .A1(\U1/aes_core/SB0/n914 ), .B0(\U1/aes_core/SB0/n868 ), .B1(
        \U1/aes_core/SB0/n1059 ), .C0(\U1/aes_core/SB0/n948 ), .C1(
        \U1/aes_core/SB0/n870 ), .Y(\U1/aes_core/SB0/n1233 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U932  ( .A0(\U1/aes_core/SB0/n1048 ), 
        .A1(\U1/aes_core/SB0/n865 ), .B0(\U1/aes_core/SB0/n845 ), .B1(
        \U1/aes_core/SB0/n844 ), .Y(\U1/aes_core/SB0/n1235 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U931  ( .A0(\U1/aes_core/SB0/n971 ), 
        .A1(\U1/aes_core/SB0/n1160 ), .B0(\U1/aes_core/SB0/n915 ), .B1(
        \U1/aes_core/SB0/n892 ), .C0(\U1/aes_core/SB0/n1235 ), .Y(
        \U1/aes_core/SB0/n1234 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U930  ( .AN(\U1/aes_core/SB0/n1231 ), 
        .B(\U1/aes_core/SB0/n1232 ), .C(\U1/aes_core/SB0/n1233 ), .D(
        \U1/aes_core/SB0/n1234 ), .Y(\U1/aes_core/SB0/n1166 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U929  ( .A(\U1/aes_core/SB0/n844 ), .B(
        \U1/aes_core/SB0/n1007 ), .Y(\U1/aes_core/SB0/n1150 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U928  ( .A0(\U1/aes_core/SB0/n937 ), .A1(
        \U1/aes_core/SB0/n844 ), .B0(\U1/aes_core/SB0/n905 ), .Y(
        \U1/aes_core/SB0/n1226 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U927  ( .A(\U1/aes_core/SB0/n905 ), .B(
        \U1/aes_core/SB0/n917 ), .Y(\U1/aes_core/SB0/n1066 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB0/U926  ( .A0(\U1/aes_core/SB0/n916 ), .A1(
        \U1/aes_core/SB0/n1160 ), .B0(\U1/aes_core/SB0/n1066 ), .B1(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1227 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U925  ( .A0(\U1/aes_core/SB0/n883 ), 
        .A1(\U1/aes_core/SB0/n843 ), .B0(\U1/aes_core/SB0/n1144 ), .B1(
        \U1/aes_core/SB0/n1051 ), .C0(\U1/aes_core/SB0/n881 ), .C1(
        \U1/aes_core/SB0/n852 ), .Y(\U1/aes_core/SB0/n1228 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U924  ( .A(\U1/aes_core/SB0/n1048 ), .Y(
        \U1/aes_core/SB0/n954 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U923  ( .A(\U1/aes_core/SB0/n850 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n928 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U922  ( .A(\U1/aes_core/SB0/n955 ), .B(
        \U1/aes_core/SB0/n1160 ), .Y(\U1/aes_core/SB0/n1127 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U921  ( .A(\U1/aes_core/SB0/n1145 ), .B(
        \U1/aes_core/SB0/n912 ), .Y(\U1/aes_core/SB0/n1107 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U920  ( .A(\U1/aes_core/SB0/n955 ), .B(
        \U1/aes_core/SB0/n914 ), .Y(\U1/aes_core/SB0/n982 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U919  ( .A(\U1/aes_core/SB0/n928 ), .B(
        \U1/aes_core/SB0/n1127 ), .C(\U1/aes_core/SB0/n1107 ), .D(
        \U1/aes_core/SB0/n982 ), .Y(\U1/aes_core/SB0/n1229 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U918  ( .A(\U1/aes_core/SB0/n935 ), .B(
        \U1/aes_core/SB0/n1048 ), .Y(\U1/aes_core/SB0/n1085 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U917  ( .A(\U1/aes_core/SB0/n949 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n1075 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U916  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n1059 ), .Y(\U1/aes_core/SB0/n1044 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U915  ( .AN(\U1/aes_core/SB0/n1085 ), 
        .B(\U1/aes_core/SB0/n1075 ), .C(\U1/aes_core/SB0/n1044 ), .Y(
        \U1/aes_core/SB0/n1230 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U914  ( .A(\U1/aes_core/SB0/n1150 ), .B(
        \U1/aes_core/SB0/n1226 ), .C(\U1/aes_core/SB0/n1227 ), .D(
        \U1/aes_core/SB0/n1228 ), .E(\U1/aes_core/SB0/n1229 ), .F(
        \U1/aes_core/SB0/n1230 ), .Y(\U1/aes_core/SB0/n837 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U913  ( .A0(\U1/aes_core/SB0/n1145 ), 
        .A1(\U1/aes_core/SB0/n891 ), .B0(\U1/aes_core/SB0/n860 ), .Y(
        \U1/aes_core/SB0/n1225 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U912  ( .A(\U1/aes_core/SB0/n1160 ), .B(
        \U1/aes_core/SB0/n1059 ), .Y(\U1/aes_core/SB0/n996 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U911  ( .A(\U1/aes_core/SB0/n916 ), .B(
        \U1/aes_core/SB0/n868 ), .Y(\U1/aes_core/SB0/n1130 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U910  ( .A(\U1/aes_core/SB0/n868 ), .B(
        \U1/aes_core/SB0/n912 ), .Y(\U1/aes_core/SB0/n1079 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U909  ( .A(\U1/aes_core/SB0/n1225 ), .B(
        \U1/aes_core/SB0/n996 ), .C(\U1/aes_core/SB0/n1130 ), .D(
        \U1/aes_core/SB0/n1079 ), .Y(\U1/aes_core/SB0/n1221 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U908  ( .A0(\U1/aes_core/SB0/n865 ), 
        .A1(\U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n1144 ), .B1(
        \U1/aes_core/SB0/n893 ), .C0(\U1/aes_core/SB0/n864 ), .C1(
        \U1/aes_core/SB0/n1007 ), .Y(\U1/aes_core/SB0/n1222 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U907  ( .A(\U1/aes_core/SB0/n913 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1098 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U906  ( .A(\U1/aes_core/SB0/n914 ), .B(
        \U1/aes_core/SB0/n862 ), .Y(\U1/aes_core/SB0/n932 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U905  ( .A(\U1/aes_core/SB0/n914 ), .B(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n1111 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U904  ( .A(\U1/aes_core/SB0/n859 ), .B(
        \U1/aes_core/SB0/n869 ), .Y(\U1/aes_core/SB0/n1149 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U903  ( .A(\U1/aes_core/SB0/n1098 ), .B(
        \U1/aes_core/SB0/n932 ), .C(\U1/aes_core/SB0/n1111 ), .D(
        \U1/aes_core/SB0/n1149 ), .Y(\U1/aes_core/SB0/n1223 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U902  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1010 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U901  ( .A(\U1/aes_core/SB0/n850 ), .B(
        \U1/aes_core/SB0/n889 ), .Y(\U1/aes_core/SB0/n1063 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U900  ( .A(\U1/aes_core/SB0/n860 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n986 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U899  ( .A(\U1/aes_core/SB0/n1133 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1163 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U898  ( .A(\U1/aes_core/SB0/n1010 ), .B(
        \U1/aes_core/SB0/n1063 ), .C(\U1/aes_core/SB0/n986 ), .D(
        \U1/aes_core/SB0/n1163 ), .Y(\U1/aes_core/SB0/n1224 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U897  ( .A(\U1/aes_core/SB0/n1221 ), .B(
        \U1/aes_core/SB0/n1222 ), .C(\U1/aes_core/SB0/n1223 ), .D(
        \U1/aes_core/SB0/n1224 ), .Y(\U1/aes_core/SB0/n1177 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U896  ( .A(\U1/aes_core/SB0/n1185 ), .B(
        \U1/aes_core/SB0/n1166 ), .C(\U1/aes_core/SB0/n837 ), .D(
        \U1/aes_core/SB0/n1177 ), .Y(\U1/aes_core/SB0/n1211 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U895  ( .A(\U1/aes_core/SB0/n883 ), .Y(
        \U1/aes_core/SB0/n959 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U894  ( .A0(\U1/aes_core/SB0/n1007 ), 
        .A1(\U1/aes_core/SB0/n1204 ), .B0(\U1/aes_core/SB0/n1064 ), .B1(
        \U1/aes_core/SB0/n852 ), .Y(\U1/aes_core/SB0/n1220 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U893  ( .A0(\U1/aes_core/SB0/n959 ), 
        .A1(\U1/aes_core/SB0/n907 ), .B0(\U1/aes_core/SB0/n858 ), .B1(
        \U1/aes_core/SB0/n850 ), .C0(\U1/aes_core/SB0/n1220 ), .Y(
        \U1/aes_core/SB0/n1212 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U892  ( .A(\U1/aes_core/SB0/n938 ), .B(
        \U1/aes_core/SB0/n935 ), .Y(\U1/aes_core/SB0/n939 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U891  ( .A0(\U1/aes_core/SB0/n1004 ), 
        .A1(\U1/aes_core/SB0/n935 ), .B0(\U1/aes_core/SB0/n1048 ), .B1(
        \U1/aes_core/SB0/n894 ), .Y(\U1/aes_core/SB0/n1219 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U890  ( .A0(\U1/aes_core/SB0/n1133 ), 
        .A1(\U1/aes_core/SB0/n939 ), .B0(\U1/aes_core/SB0/n888 ), .B1(
        \U1/aes_core/SB0/n869 ), .C0(\U1/aes_core/SB0/n1219 ), .Y(
        \U1/aes_core/SB0/n1213 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U889  ( .A(\U1/aes_core/SB0/n864 ), .B(
        \U1/aes_core/SB0/n1005 ), .Y(\U1/aes_core/SB0/n1215 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U888  ( .A(\U1/aes_core/SB0/n914 ), .B(
        \U1/aes_core/SB0/n889 ), .Y(\U1/aes_core/SB0/n947 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U887  ( .A(\U1/aes_core/SB0/n947 ), .Y(
        \U1/aes_core/SB0/n1216 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U886  ( .A(\U1/aes_core/SB0/n956 ), .B(
        \U1/aes_core/SB0/n883 ), .Y(\U1/aes_core/SB0/n1101 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U885  ( .A(\U1/aes_core/SB0/n878 ), .B(
        \U1/aes_core/SB0/n880 ), .Y(\U1/aes_core/SB0/n922 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U883  ( .A(\U1/aes_core/SB0/n907 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n1091 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U881  ( .A0(\U1/aes_core/SB0/n948 ), 
        .A1(\U1/aes_core/SB0/n1215 ), .B0(\U1/aes_core/SB0/n971 ), .B1(
        \U1/aes_core/SB0/n1216 ), .C0(\U1/aes_core/SB0/n1217 ), .Y(
        \U1/aes_core/SB0/n1214 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U880  ( .AN(\U1/aes_core/SB0/n1211 ), 
        .B(\U1/aes_core/SB0/n1212 ), .C(\U1/aes_core/SB0/n1213 ), .D(
        \U1/aes_core/SB0/n1214 ), .Y(\U1/aes_core/sb0 [16]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U879  ( .A(\U1/aes_core/SB0/n935 ), .B(
        \U1/aes_core/SB0/n1144 ), .Y(\U1/aes_core/SB0/n1084 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U878  ( .A(\U1/aes_core/SB0/n988 ), .B(
        \U1/aes_core/SB0/n938 ), .Y(\U1/aes_core/SB0/n1124 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U877  ( .A(\U1/aes_core/SB0/n971 ), .B(
        \U1/aes_core/SB0/n860 ), .Y(\U1/aes_core/SB0/n989 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U876  ( .A0(\U1/aes_core/SB0/n989 ), .A1(
        \U1/aes_core/SB0/n935 ), .B0(\U1/aes_core/SB0/n846 ), .Y(
        \U1/aes_core/SB0/n1206 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U875  ( .A(\U1/aes_core/SB0/n907 ), .B(
        \U1/aes_core/SB0/n859 ), .Y(\U1/aes_core/SB0/n1108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U874  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n907 ), .Y(\U1/aes_core/SB0/n983 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U873  ( .A(\U1/aes_core/SB0/n862 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n1076 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U872  ( .A(\U1/aes_core/SB0/n1108 ), .B(
        \U1/aes_core/SB0/n983 ), .C(\U1/aes_core/SB0/n1076 ), .Y(
        \U1/aes_core/SB0/n1207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U871  ( .A(\U1/aes_core/SB0/n907 ), .B(
        \U1/aes_core/SB0/n848 ), .Y(\U1/aes_core/SB0/n1049 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U870  ( .A(\U1/aes_core/SB0/n862 ), .B(
        \U1/aes_core/SB0/n871 ), .C(\U1/aes_core/SB0/n850 ), .Y(
        \U1/aes_core/SB0/n1210 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U869  ( .A0(\U1/aes_core/SB0/n1049 ), 
        .A1(\U1/aes_core/SB0/n882 ), .B0(\U1/aes_core/SB0/n1210 ), .B1(
        \U1/aes_core/SB0/n852 ), .C0(\U1/aes_core/SB0/n988 ), .C1(
        \U1/aes_core/SB0/n956 ), .Y(\U1/aes_core/SB0/n1208 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U868  ( .A0(\U1/aes_core/SB0/n881 ), .A1(
        \U1/aes_core/SB0/n853 ), .B0(\U1/aes_core/SB0/n880 ), .B1(
        \U1/aes_core/SB0/n883 ), .Y(\U1/aes_core/SB0/n1209 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U867  ( .A(\U1/aes_core/SB0/n1084 ), .B(
        \U1/aes_core/SB0/n1124 ), .C(\U1/aes_core/SB0/n1206 ), .D(
        \U1/aes_core/SB0/n1207 ), .E(\U1/aes_core/SB0/n1208 ), .F(
        \U1/aes_core/SB0/n1209 ), .Y(\U1/aes_core/SB0/n838 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U866  ( .A(\U1/aes_core/SB0/n1007 ), .B(
        \U1/aes_core/SB0/n1048 ), .Y(\U1/aes_core/SB0/n1159 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U865  ( .A0(\U1/aes_core/SB0/n1007 ), 
        .A1(\U1/aes_core/SB0/n917 ), .B0(\U1/aes_core/SB0/n1144 ), .Y(
        \U1/aes_core/SB0/n1198 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U864  ( .A(\U1/aes_core/SB0/n913 ), .B(
        \U1/aes_core/SB0/n907 ), .Y(\U1/aes_core/SB0/n1156 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U863  ( .A0(\U1/aes_core/SB0/n1051 ), 
        .A1(\U1/aes_core/SB0/n878 ), .B0(\U1/aes_core/SB0/n1156 ), .B1(
        \U1/aes_core/SB0/n864 ), .Y(\U1/aes_core/SB0/n1199 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U862  ( .A0(\U1/aes_core/SB0/n1064 ), 
        .A1(\U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n894 ), .B1(
        \U1/aes_core/SB0/n988 ), .C0(\U1/aes_core/SB0/n880 ), .C1(
        \U1/aes_core/SB0/n937 ), .Y(\U1/aes_core/SB0/n1200 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U861  ( .A(\U1/aes_core/SB0/n845 ), .B(
        \U1/aes_core/SB0/n1205 ), .Y(\U1/aes_core/SB0/n1100 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U860  ( .A(\U1/aes_core/SB0/n858 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1093 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U859  ( .A(\U1/aes_core/SB0/n916 ), .B(
        \U1/aes_core/SB0/n863 ), .Y(\U1/aes_core/SB0/n1083 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U858  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n848 ), .Y(\U1/aes_core/SB0/n953 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U857  ( .AN(\U1/aes_core/SB0/n1100 ), 
        .B(\U1/aes_core/SB0/n1093 ), .C(\U1/aes_core/SB0/n1083 ), .D(
        \U1/aes_core/SB0/n953 ), .Y(\U1/aes_core/SB0/n1201 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U856  ( .A(\U1/aes_core/SB0/n956 ), .B(
        \U1/aes_core/SB0/n1204 ), .Y(\U1/aes_core/SB0/n974 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U855  ( .A(\U1/aes_core/SB0/n878 ), .B(
        \U1/aes_core/SB0/n894 ), .Y(\U1/aes_core/SB0/n921 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U853  ( .A(\U1/aes_core/SB0/n1160 ), .B(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n1134 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U851  ( .A(\U1/aes_core/SB0/n1159 ), .B(
        \U1/aes_core/SB0/n1198 ), .C(\U1/aes_core/SB0/n1199 ), .D(
        \U1/aes_core/SB0/n1200 ), .E(\U1/aes_core/SB0/n1201 ), .F(
        \U1/aes_core/SB0/n1202 ), .Y(\U1/aes_core/SB0/n1165 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U850  ( .A(\U1/aes_core/SB0/n940 ), .B(
        \U1/aes_core/SB0/n1144 ), .Y(\U1/aes_core/SB0/n1146 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U849  ( .A(\U1/aes_core/SB0/n988 ), .B(
        \U1/aes_core/SB0/n1064 ), .Y(\U1/aes_core/SB0/n908 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U848  ( .A(\U1/aes_core/SB0/n1007 ), .B(
        \U1/aes_core/SB0/n937 ), .Y(\U1/aes_core/SB0/n1096 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U847  ( .A(\U1/aes_core/SB0/n843 ), .B(
        \U1/aes_core/SB0/n937 ), .Y(\U1/aes_core/SB0/n1081 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U846  ( .A(\U1/aes_core/SB0/n912 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n995 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U845  ( .A(\U1/aes_core/SB0/n862 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1129 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U844  ( .A(\U1/aes_core/SB0/n858 ), .B(
        \U1/aes_core/SB0/n862 ), .Y(\U1/aes_core/SB0/n1009 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U843  ( .A(\U1/aes_core/SB0/n948 ), .B(
        \U1/aes_core/SB0/n891 ), .Y(\U1/aes_core/SB0/n1110 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U842  ( .A(\U1/aes_core/SB0/n995 ), .B(
        \U1/aes_core/SB0/n1129 ), .C(\U1/aes_core/SB0/n1009 ), .D(
        \U1/aes_core/SB0/n1110 ), .Y(\U1/aes_core/SB0/n1194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U841  ( .A(\U1/aes_core/SB0/n843 ), .B(
        \U1/aes_core/SB0/n1048 ), .Y(\U1/aes_core/SB0/n1060 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U840  ( .A(\U1/aes_core/SB0/n844 ), .B(
        \U1/aes_core/SB0/n1064 ), .Y(\U1/aes_core/SB0/n934 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U839  ( .A(\U1/aes_core/SB0/n917 ), .B(
        \U1/aes_core/SB0/n878 ), .Y(\U1/aes_core/SB0/n984 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U838  ( .A(\U1/aes_core/SB0/n956 ), .B(
        \U1/aes_core/SB0/n878 ), .Y(\U1/aes_core/SB0/n1161 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U837  ( .A0(\U1/aes_core/SB0/n878 ), .A1(
        \U1/aes_core/SB0/n843 ), .B0(\U1/aes_core/SB0/n1048 ), .B1(
        \U1/aes_core/SB0/n917 ), .Y(\U1/aes_core/SB0/n1196 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U836  ( .A0(\U1/aes_core/SB0/n1064 ), 
        .A1(\U1/aes_core/SB0/n846 ), .B0(\U1/aes_core/SB0/n1051 ), .B1(
        \U1/aes_core/SB0/n988 ), .Y(\U1/aes_core/SB0/n1197 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U835  ( .A(\U1/aes_core/SB0/n1060 ), .B(
        \U1/aes_core/SB0/n934 ), .C(\U1/aes_core/SB0/n984 ), .D(
        \U1/aes_core/SB0/n1161 ), .E(\U1/aes_core/SB0/n1196 ), .F(
        \U1/aes_core/SB0/n1197 ), .Y(\U1/aes_core/SB0/n1195 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U834  ( .A(\U1/aes_core/SB0/n1146 ), .B(
        \U1/aes_core/SB0/n908 ), .C(\U1/aes_core/SB0/n1096 ), .D(
        \U1/aes_core/SB0/n1081 ), .E(\U1/aes_core/SB0/n1194 ), .F(
        \U1/aes_core/SB0/n1195 ), .Y(\U1/aes_core/SB0/n1176 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U833  ( .A0(\U1/aes_core/SB0/n912 ), 
        .A1(\U1/aes_core/SB0/n915 ), .B0(\U1/aes_core/SB0/n859 ), .B1(
        \U1/aes_core/SB0/n971 ), .C0(\U1/aes_core/SB0/n1176 ), .Y(
        \U1/aes_core/SB0/n1193 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U832  ( .A(\U1/aes_core/SB0/n1193 ), .Y(
        \U1/aes_core/SB0/n1186 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U831  ( .A(\U1/aes_core/SB0/n880 ), .B(
        \U1/aes_core/SB0/n917 ), .Y(\U1/aes_core/SB0/n890 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U830  ( .A0(\U1/aes_core/SB0/n913 ), .A1(
        \U1/aes_core/SB0/n890 ), .B0(\U1/aes_core/SB0/n858 ), .Y(
        \U1/aes_core/SB0/n1190 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U829  ( .A0(\U1/aes_core/SB0/n948 ), .A1(
        \U1/aes_core/SB0/n869 ), .B0(\U1/aes_core/SB0/n906 ), .Y(
        \U1/aes_core/SB0/n1191 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U828  ( .A0(\U1/aes_core/SB0/n949 ), .A1(
        \U1/aes_core/SB0/n907 ), .B0(\U1/aes_core/SB0/n863 ), .Y(
        \U1/aes_core/SB0/n1192 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U827  ( .A(\U1/aes_core/SB0/n916 ), .B(
        \U1/aes_core/SB0/n870 ), .Y(\U1/aes_core/SB0/n1117 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U826  ( .A(\U1/aes_core/SB0/n1190 ), .B(
        \U1/aes_core/SB0/n1191 ), .C(\U1/aes_core/SB0/n1192 ), .D(
        \U1/aes_core/SB0/n1117 ), .Y(\U1/aes_core/SB0/n1187 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U825  ( .A(\U1/aes_core/SB0/n871 ), .B(
        \U1/aes_core/SB0/n955 ), .Y(\U1/aes_core/SB0/n901 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB0/U824  ( .A(\U1/aes_core/SB0/n901 ), .B(
        \U1/aes_core/SB0/n881 ), .C(\U1/aes_core/SB0/n894 ), .Y(
        \U1/aes_core/SB0/n1189 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U823  ( .A0(\U1/aes_core/SB0/n917 ), 
        .A1(\U1/aes_core/SB0/n844 ), .B0(\U1/aes_core/SB0/n1189 ), .B1(
        \U1/aes_core/SB0/n883 ), .C0(\U1/aes_core/SB0/n845 ), .C1(
        \U1/aes_core/SB0/n853 ), .Y(\U1/aes_core/SB0/n1188 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U822  ( .A(\U1/aes_core/SB0/n838 ), .B(
        \U1/aes_core/SB0/n1165 ), .C(\U1/aes_core/SB0/n1185 ), .D(
        \U1/aes_core/SB0/n1186 ), .E(\U1/aes_core/SB0/n1187 ), .F(
        \U1/aes_core/SB0/n1188 ), .Y(\U1/aes_core/sb0 [17]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U821  ( .A0(\U1/aes_core/SB0/n889 ), .A1(
        \U1/aes_core/SB0/n869 ), .B0(\U1/aes_core/SB0/n848 ), .B1(
        \U1/aes_core/SB0/n858 ), .Y(\U1/aes_core/SB0/n1184 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U820  ( .A0(\U1/aes_core/SB0/n938 ), 
        .A1(\U1/aes_core/SB0/n844 ), .B0(\U1/aes_core/SB0/n988 ), .B1(
        \U1/aes_core/SB0/n917 ), .C0(\U1/aes_core/SB0/n1184 ), .Y(
        \U1/aes_core/SB0/n1178 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U819  ( .A(\U1/aes_core/SB0/n863 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1080 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U818  ( .A(\U1/aes_core/SB0/n889 ), .B(
        \U1/aes_core/SB0/n913 ), .Y(\U1/aes_core/SB0/n1099 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U817  ( .A(\U1/aes_core/SB0/n869 ), .B(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n1131 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U816  ( .A(\U1/aes_core/SB0/n949 ), .B(
        \U1/aes_core/SB0/n906 ), .Y(\U1/aes_core/SB0/n1112 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U815  ( .A(\U1/aes_core/SB0/n1080 ), .B(
        \U1/aes_core/SB0/n1099 ), .C(\U1/aes_core/SB0/n1131 ), .D(
        \U1/aes_core/SB0/n1112 ), .Y(\U1/aes_core/SB0/n1179 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U814  ( .A(\U1/aes_core/SB0/n843 ), .B(
        \U1/aes_core/SB0/n865 ), .Y(\U1/aes_core/SB0/n960 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U813  ( .A0(\U1/aes_core/SB0/n912 ), .A1(
        \U1/aes_core/SB0/n960 ), .B0(\U1/aes_core/SB0/n859 ), .Y(
        \U1/aes_core/SB0/n1181 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U812  ( .A0(\U1/aes_core/SB0/n862 ), .A1(
        \U1/aes_core/SB0/n971 ), .B0(\U1/aes_core/SB0/n959 ), .Y(
        \U1/aes_core/SB0/n1182 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U811  ( .A0(\U1/aes_core/SB0/n954 ), .A1(
        \U1/aes_core/SB0/n914 ), .B0(\U1/aes_core/SB0/n860 ), .Y(
        \U1/aes_core/SB0/n1183 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U810  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n862 ), .Y(\U1/aes_core/SB0/n987 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U809  ( .A(\U1/aes_core/SB0/n1181 ), .B(
        \U1/aes_core/SB0/n1182 ), .C(\U1/aes_core/SB0/n1183 ), .D(
        \U1/aes_core/SB0/n987 ), .Y(\U1/aes_core/SB0/n1180 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U808  ( .A(\U1/aes_core/SB0/n1175 ), .B(
        \U1/aes_core/SB0/n1176 ), .C(\U1/aes_core/SB0/n1177 ), .D(
        \U1/aes_core/SB0/n1178 ), .E(\U1/aes_core/SB0/n1179 ), .F(
        \U1/aes_core/SB0/n1180 ), .Y(\U1/aes_core/SB0/n839 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U807  ( .A0(\U1/aes_core/SB0/n1059 ), 
        .A1(\U1/aes_core/SB0/n858 ), .B0(\U1/aes_core/SB0/n850 ), .B1(
        \U1/aes_core/SB0/n915 ), .C0(\U1/aes_core/SB0/n839 ), .Y(
        \U1/aes_core/SB0/n1174 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U806  ( .A(\U1/aes_core/SB0/n1174 ), .Y(
        \U1/aes_core/SB0/n1167 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U805  ( .A(\U1/aes_core/SB0/n906 ), .B(
        \U1/aes_core/SB0/n1145 ), .Y(\U1/aes_core/SB0/n997 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U804  ( .A1N(\U1/aes_core/SB0/n997 ), 
        .A0(\U1/aes_core/SB0/n888 ), .B0(\U1/aes_core/SB0/n916 ), .Y(
        \U1/aes_core/SB0/n1171 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U803  ( .A0(\U1/aes_core/SB0/n948 ), .A1(
        \U1/aes_core/SB0/n1066 ), .B0(\U1/aes_core/SB0/n889 ), .Y(
        \U1/aes_core/SB0/n1172 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U802  ( .A0(\U1/aes_core/SB0/n862 ), .A1(
        \U1/aes_core/SB0/n907 ), .B0(\U1/aes_core/SB0/n868 ), .Y(
        \U1/aes_core/SB0/n1173 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U801  ( .A(\U1/aes_core/SB0/n891 ), .B(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n1116 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U800  ( .A(\U1/aes_core/SB0/n1171 ), .B(
        \U1/aes_core/SB0/n1172 ), .C(\U1/aes_core/SB0/n1173 ), .D(
        \U1/aes_core/SB0/n1116 ), .Y(\U1/aes_core/SB0/n1168 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U799  ( .A(\U1/aes_core/SB0/n892 ), .B(
        \U1/aes_core/SB0/n860 ), .Y(\U1/aes_core/SB0/n861 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U798  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n914 ), .Y(\U1/aes_core/SB0/n1170 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U797  ( .A0(\U1/aes_core/SB0/n861 ), 
        .A1(\U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n1170 ), .B1(
        \U1/aes_core/SB0/n880 ), .C0(\U1/aes_core/SB0/n937 ), .C1(
        \U1/aes_core/SB0/n935 ), .Y(\U1/aes_core/SB0/n1169 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U796  ( .A(\U1/aes_core/SB0/n1164 ), .B(
        \U1/aes_core/SB0/n1165 ), .C(\U1/aes_core/SB0/n1166 ), .D(
        \U1/aes_core/SB0/n1167 ), .E(\U1/aes_core/SB0/n1168 ), .F(
        \U1/aes_core/SB0/n1169 ), .Y(\U1/aes_core/sb0 [18]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U795  ( .A(\U1/aes_core/SB0/n1059 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n856 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U794  ( .AN(\U1/aes_core/SB0/n1161 ), 
        .B(\U1/aes_core/SB0/n1162 ), .C(\U1/aes_core/SB0/n1163 ), .D(
        \U1/aes_core/SB0/n856 ), .Y(\U1/aes_core/SB0/n1153 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U793  ( .A0(\U1/aes_core/SB0/n1160 ), 
        .A1(\U1/aes_core/SB0/n889 ), .B0(\U1/aes_core/SB0/n971 ), .Y(
        \U1/aes_core/SB0/n1157 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U790  ( .A(\U1/aes_core/SB0/n915 ), .B(
        \U1/aes_core/SB0/n868 ), .Y(\U1/aes_core/SB0/n904 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U789  ( .A0(\U1/aes_core/SB0/n1051 ), 
        .A1(\U1/aes_core/SB0/n846 ), .B0(\U1/aes_core/SB0/n904 ), .B1(
        \U1/aes_core/SB0/n893 ), .C0(\U1/aes_core/SB0/n852 ), .C1(
        \U1/aes_core/SB0/n843 ), .Y(\U1/aes_core/SB0/n1155 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U788  ( .A(\U1/aes_core/SB0/n1150 ), .B(
        \U1/aes_core/SB0/n1151 ), .C(\U1/aes_core/SB0/n1152 ), .D(
        \U1/aes_core/SB0/n1153 ), .E(\U1/aes_core/SB0/n1154 ), .F(
        \U1/aes_core/SB0/n1155 ), .Y(\U1/aes_core/SB0/n941 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U787  ( .AN(\U1/aes_core/SB0/n1146 ), 
        .B(\U1/aes_core/SB0/n1147 ), .C(\U1/aes_core/SB0/n1148 ), .D(
        \U1/aes_core/SB0/n1149 ), .Y(\U1/aes_core/SB0/n1136 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U786  ( .A0(\U1/aes_core/SB0/n858 ), 
        .A1(\U1/aes_core/SB0/n948 ), .B0(\U1/aes_core/SB0/n863 ), .B1(
        \U1/aes_core/SB0/n949 ), .C0(\U1/aes_core/SB0/n1145 ), .C1(
        \U1/aes_core/SB0/n848 ), .Y(\U1/aes_core/SB0/n1137 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U785  ( .A0(\U1/aes_core/SB0/n894 ), .A1(
        \U1/aes_core/SB0/n988 ), .B0(\U1/aes_core/SB0/n1144 ), .B1(
        \U1/aes_core/SB0/n1051 ), .Y(\U1/aes_core/SB0/n1143 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U784  ( .A0(\U1/aes_core/SB0/n971 ), 
        .A1(\U1/aes_core/SB0/n954 ), .B0(\U1/aes_core/SB0/n955 ), .B1(
        \U1/aes_core/SB0/n891 ), .C0(\U1/aes_core/SB0/n1143 ), .Y(
        \U1/aes_core/SB0/n1138 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U783  ( .A(\U1/aes_core/SB0/n883 ), .B(
        \U1/aes_core/SB0/n844 ), .Y(\U1/aes_core/SB0/n1141 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U782  ( .A0(\U1/aes_core/SB0/n1059 ), 
        .A1(\U1/aes_core/SB0/n1140 ), .B0(\U1/aes_core/SB0/n862 ), .B1(
        \U1/aes_core/SB0/n1141 ), .C0(\U1/aes_core/SB0/n1142 ), .Y(
        \U1/aes_core/SB0/n1139 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U781  ( .AN(\U1/aes_core/SB0/n1136 ), 
        .B(\U1/aes_core/SB0/n1137 ), .C(\U1/aes_core/SB0/n1138 ), .D(
        \U1/aes_core/SB0/n1139 ), .Y(\U1/aes_core/SB0/n896 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U780  ( .A(\U1/aes_core/SB0/n1135 ), .Y(
        \U1/aes_core/SB0/n1119 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U779  ( .A0(\U1/aes_core/SB0/n1004 ), 
        .A1(\U1/aes_core/SB0/n935 ), .B0(\U1/aes_core/SB0/n1134 ), .Y(
        \U1/aes_core/SB0/n1120 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U778  ( .A0(\U1/aes_core/SB0/n862 ), .A1(
        \U1/aes_core/SB0/n863 ), .B0(\U1/aes_core/SB0/n892 ), .B1(
        \U1/aes_core/SB0/n1133 ), .Y(\U1/aes_core/SB0/n1132 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U777  ( .A0(\U1/aes_core/SB0/n881 ), 
        .A1(\U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n865 ), .B1(
        \U1/aes_core/SB0/n853 ), .C0(\U1/aes_core/SB0/n1132 ), .Y(
        \U1/aes_core/SB0/n1121 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U776  ( .A(\U1/aes_core/SB0/n1128 ), .B(
        \U1/aes_core/SB0/n1129 ), .C(\U1/aes_core/SB0/n1130 ), .D(
        \U1/aes_core/SB0/n1131 ), .Y(\U1/aes_core/SB0/n1122 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U775  ( .AN(\U1/aes_core/SB0/n1124 ), 
        .B(\U1/aes_core/SB0/n1125 ), .C(\U1/aes_core/SB0/n1126 ), .D(
        \U1/aes_core/SB0/n1127 ), .Y(\U1/aes_core/SB0/n1123 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U774  ( .A(\U1/aes_core/SB0/n1118 ), .B(
        \U1/aes_core/SB0/n1119 ), .C(\U1/aes_core/SB0/n1120 ), .D(
        \U1/aes_core/SB0/n1121 ), .E(\U1/aes_core/SB0/n1122 ), .F(
        \U1/aes_core/SB0/n1123 ), .Y(\U1/aes_core/SB0/n992 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U773  ( .A0(\U1/aes_core/SB0/n905 ), .A1(
        \U1/aes_core/SB0/n988 ), .B0(\U1/aes_core/SB0/n1117 ), .Y(
        \U1/aes_core/SB0/n1102 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U772  ( .AN(\U1/aes_core/SB0/n1113 ), 
        .B(\U1/aes_core/SB0/n1114 ), .C(\U1/aes_core/SB0/n1115 ), .D(
        \U1/aes_core/SB0/n1116 ), .Y(\U1/aes_core/SB0/n1103 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U771  ( .A(\U1/aes_core/SB0/n871 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n857 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U770  ( .A(\U1/aes_core/SB0/n1110 ), .B(
        \U1/aes_core/SB0/n1111 ), .C(\U1/aes_core/SB0/n1112 ), .D(
        \U1/aes_core/SB0/n857 ), .Y(\U1/aes_core/SB0/n1104 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U769  ( .A(\U1/aes_core/SB0/n1106 ), .B(
        \U1/aes_core/SB0/n1107 ), .C(\U1/aes_core/SB0/n1108 ), .D(
        \U1/aes_core/SB0/n1109 ), .Y(\U1/aes_core/SB0/n1105 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U768  ( .A(\U1/aes_core/SB0/n1100 ), .B(
        \U1/aes_core/SB0/n1101 ), .C(\U1/aes_core/SB0/n1102 ), .D(
        \U1/aes_core/SB0/n1103 ), .E(\U1/aes_core/SB0/n1104 ), .F(
        \U1/aes_core/SB0/n1105 ), .Y(\U1/aes_core/SB0/n968 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U767  ( .AN(\U1/aes_core/SB0/n1096 ), 
        .B(\U1/aes_core/SB0/n1097 ), .C(\U1/aes_core/SB0/n1098 ), .D(
        \U1/aes_core/SB0/n1099 ), .Y(\U1/aes_core/SB0/n1087 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U766  ( .A(\U1/aes_core/SB0/n1092 ), .B(
        \U1/aes_core/SB0/n1093 ), .C(\U1/aes_core/SB0/n1094 ), .D(
        \U1/aes_core/SB0/n1095 ), .Y(\U1/aes_core/SB0/n1088 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U765  ( .A(\U1/aes_core/SB0/n906 ), .B(
        \U1/aes_core/SB0/n870 ), .C(\U1/aes_core/SB0/n868 ), .Y(
        \U1/aes_core/SB0/n1090 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U764  ( .A0(\U1/aes_core/SB0/n1090 ), 
        .A1(\U1/aes_core/SB0/n880 ), .B0(\U1/aes_core/SB0/n1051 ), .B1(
        \U1/aes_core/SB0/n844 ), .C0(\U1/aes_core/SB0/n1091 ), .Y(
        \U1/aes_core/SB0/n1089 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U763  ( .A(\U1/aes_core/SB0/n1084 ), .B(
        \U1/aes_core/SB0/n1085 ), .C(\U1/aes_core/SB0/n1086 ), .D(
        \U1/aes_core/SB0/n1087 ), .E(\U1/aes_core/SB0/n1088 ), .F(
        \U1/aes_core/SB0/n1089 ), .Y(\U1/aes_core/SB0/n920 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U762  ( .A0(\U1/aes_core/SB0/n1051 ), 
        .A1(\U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n1083 ), .Y(
        \U1/aes_core/SB0/n1069 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U761  ( .A0(\U1/aes_core/SB0/n916 ), .A1(
        \U1/aes_core/SB0/n914 ), .B0(\U1/aes_core/SB0/n859 ), .B1(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n1082 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U760  ( .A0(\U1/aes_core/SB0/n1005 ), 
        .A1(\U1/aes_core/SB0/n917 ), .B0(\U1/aes_core/SB0/n1004 ), .B1(
        \U1/aes_core/SB0/n940 ), .C0(\U1/aes_core/SB0/n1082 ), .Y(
        \U1/aes_core/SB0/n1070 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U759  ( .A(\U1/aes_core/SB0/n1081 ), .Y(
        \U1/aes_core/SB0/n1078 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U758  ( .AN(\U1/aes_core/SB0/n1077 ), 
        .B(\U1/aes_core/SB0/n1078 ), .C(\U1/aes_core/SB0/n1079 ), .D(
        \U1/aes_core/SB0/n1080 ), .Y(\U1/aes_core/SB0/n1071 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U757  ( .A(\U1/aes_core/SB0/n1073 ), .B(
        \U1/aes_core/SB0/n1074 ), .C(\U1/aes_core/SB0/n1075 ), .D(
        \U1/aes_core/SB0/n1076 ), .Y(\U1/aes_core/SB0/n1072 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U756  ( .A(\U1/aes_core/SB0/n1067 ), .B(
        \U1/aes_core/SB0/n1068 ), .C(\U1/aes_core/SB0/n1069 ), .D(
        \U1/aes_core/SB0/n1070 ), .E(\U1/aes_core/SB0/n1071 ), .F(
        \U1/aes_core/SB0/n1072 ), .Y(\U1/aes_core/SB0/n961 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U755  ( .A0(\U1/aes_core/SB0/n870 ), .A1(
        \U1/aes_core/SB0/n1066 ), .B0(\U1/aes_core/SB0/n860 ), .B1(
        \U1/aes_core/SB0/n914 ), .Y(\U1/aes_core/SB0/n1065 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U754  ( .A0(\U1/aes_core/SB0/n988 ), 
        .A1(\U1/aes_core/SB0/n843 ), .B0(\U1/aes_core/SB0/n1064 ), .B1(
        \U1/aes_core/SB0/n853 ), .C0(\U1/aes_core/SB0/n1065 ), .Y(
        \U1/aes_core/SB0/n1052 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U753  ( .AN(\U1/aes_core/SB0/n1060 ), 
        .B(\U1/aes_core/SB0/n1061 ), .C(\U1/aes_core/SB0/n1062 ), .D(
        \U1/aes_core/SB0/n1063 ), .Y(\U1/aes_core/SB0/n1053 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U752  ( .A0(\U1/aes_core/SB0/n850 ), .A1(
        \U1/aes_core/SB0/n1059 ), .B0(\U1/aes_core/SB0/n859 ), .Y(
        \U1/aes_core/SB0/n1055 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U751  ( .A(\U1/aes_core/SB0/n883 ), .B(
        \U1/aes_core/SB0/n878 ), .Y(\U1/aes_core/SB0/n1058 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U750  ( .A0(\U1/aes_core/SB0/n907 ), .A1(
        \U1/aes_core/SB0/n1058 ), .B0(\U1/aes_core/SB0/n906 ), .B1(
        \U1/aes_core/SB0/n960 ), .Y(\U1/aes_core/SB0/n1057 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U749  ( .A(\U1/aes_core/SB0/n1055 ), .B(
        \U1/aes_core/SB0/n1056 ), .C(\U1/aes_core/SB0/n1057 ), .Y(
        \U1/aes_core/SB0/n1054 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U748  ( .A(\U1/aes_core/SB0/n968 ), .B(
        \U1/aes_core/SB0/n920 ), .C(\U1/aes_core/SB0/n961 ), .D(
        \U1/aes_core/SB0/n1052 ), .E(\U1/aes_core/SB0/n1053 ), .F(
        \U1/aes_core/SB0/n1054 ), .Y(\U1/aes_core/SB0/n874 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U747  ( .A(\U1/aes_core/SB0/n941 ), .B(
        \U1/aes_core/SB0/n896 ), .C(\U1/aes_core/SB0/n992 ), .D(
        \U1/aes_core/SB0/n874 ), .Y(\U1/aes_core/SB0/n1038 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U746  ( .A0(\U1/aes_core/SB0/n894 ), .A1(
        \U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n1051 ), .B1(
        \U1/aes_core/SB0/n878 ), .Y(\U1/aes_core/SB0/n1050 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U745  ( .A0(\U1/aes_core/SB0/n889 ), 
        .A1(\U1/aes_core/SB0/n871 ), .B0(\U1/aes_core/SB0/n858 ), .B1(
        \U1/aes_core/SB0/n850 ), .C0(\U1/aes_core/SB0/n1050 ), .Y(
        \U1/aes_core/SB0/n1039 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U744  ( .A(\U1/aes_core/SB0/n1049 ), .Y(
        \U1/aes_core/SB0/n1046 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U743  ( .A0(\U1/aes_core/SB0/n1048 ), 
        .A1(\U1/aes_core/SB0/n917 ), .B0(\U1/aes_core/SB0/n989 ), .B1(
        \U1/aes_core/SB0/n937 ), .Y(\U1/aes_core/SB0/n1047 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U742  ( .A0(\U1/aes_core/SB0/n870 ), 
        .A1(\U1/aes_core/SB0/n1046 ), .B0(\U1/aes_core/SB0/n888 ), .B1(
        \U1/aes_core/SB0/n939 ), .C0(\U1/aes_core/SB0/n1047 ), .Y(
        \U1/aes_core/SB0/n1040 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U741  ( .A0(\U1/aes_core/SB0/n848 ), .A1(
        \U1/aes_core/SB0/n971 ), .B0(\U1/aes_core/SB0/n868 ), .Y(
        \U1/aes_core/SB0/n1042 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB0/U740  ( .A(\U1/aes_core/SB0/n1042 ), .B(
        \U1/aes_core/SB0/n1043 ), .C(\U1/aes_core/SB0/n1044 ), .D(
        \U1/aes_core/SB0/n1045 ), .Y(\U1/aes_core/SB0/n1041 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U739  ( .AN(\U1/aes_core/SB0/n1038 ), 
        .B(\U1/aes_core/SB0/n1039 ), .C(\U1/aes_core/SB0/n1040 ), .D(
        \U1/aes_core/SB0/n1041 ), .Y(\U1/aes_core/sb0 [19]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U738  ( .A(\U1/aes_core/SB0/n188 ), .B(
        \U1/aes_core/SB0/n371 ), .Y(\U1/aes_core/SB0/n311 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U737  ( .A(\U1/aes_core/SB0/n241 ), .B(
        \U1/aes_core/SB0/n191 ), .Y(\U1/aes_core/SB0/n351 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U736  ( .A(\U1/aes_core/SB0/n224 ), .B(
        \U1/aes_core/SB0/n113 ), .Y(\U1/aes_core/SB0/n242 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U735  ( .A0(\U1/aes_core/SB0/n242 ), .A1(
        \U1/aes_core/SB0/n188 ), .B0(\U1/aes_core/SB0/n99 ), .Y(
        \U1/aes_core/SB0/n1033 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U734  ( .A(\U1/aes_core/SB0/n160 ), .B(
        \U1/aes_core/SB0/n112 ), .Y(\U1/aes_core/SB0/n335 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U733  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n160 ), .Y(\U1/aes_core/SB0/n236 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U732  ( .A(\U1/aes_core/SB0/n115 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n303 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U731  ( .A(\U1/aes_core/SB0/n335 ), .B(
        \U1/aes_core/SB0/n236 ), .C(\U1/aes_core/SB0/n303 ), .Y(
        \U1/aes_core/SB0/n1034 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U730  ( .A(\U1/aes_core/SB0/n160 ), .B(
        \U1/aes_core/SB0/n101 ), .Y(\U1/aes_core/SB0/n276 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U729  ( .A(\U1/aes_core/SB0/n115 ), .B(
        \U1/aes_core/SB0/n124 ), .C(\U1/aes_core/SB0/n103 ), .Y(
        \U1/aes_core/SB0/n1037 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U728  ( .A0(\U1/aes_core/SB0/n276 ), 
        .A1(\U1/aes_core/SB0/n135 ), .B0(\U1/aes_core/SB0/n1037 ), .B1(
        \U1/aes_core/SB0/n105 ), .C0(\U1/aes_core/SB0/n241 ), .C1(
        \U1/aes_core/SB0/n209 ), .Y(\U1/aes_core/SB0/n1035 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U727  ( .A0(\U1/aes_core/SB0/n134 ), .A1(
        \U1/aes_core/SB0/n106 ), .B0(\U1/aes_core/SB0/n133 ), .B1(
        \U1/aes_core/SB0/n136 ), .Y(\U1/aes_core/SB0/n1036 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U726  ( .A(\U1/aes_core/SB0/n311 ), .B(
        \U1/aes_core/SB0/n351 ), .C(\U1/aes_core/SB0/n1033 ), .D(
        \U1/aes_core/SB0/n1034 ), .E(\U1/aes_core/SB0/n1035 ), .F(
        \U1/aes_core/SB0/n1036 ), .Y(\U1/aes_core/SB0/n91 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U725  ( .A(\U1/aes_core/SB0/n260 ), .B(
        \U1/aes_core/SB0/n275 ), .Y(\U1/aes_core/SB0/n386 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U724  ( .A0(\U1/aes_core/SB0/n260 ), .A1(
        \U1/aes_core/SB0/n170 ), .B0(\U1/aes_core/SB0/n371 ), .Y(
        \U1/aes_core/SB0/n1025 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U723  ( .A(\U1/aes_core/SB0/n166 ), .B(
        \U1/aes_core/SB0/n160 ), .Y(\U1/aes_core/SB0/n383 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U722  ( .A0(\U1/aes_core/SB0/n278 ), .A1(
        \U1/aes_core/SB0/n131 ), .B0(\U1/aes_core/SB0/n383 ), .B1(
        \U1/aes_core/SB0/n117 ), .Y(\U1/aes_core/SB0/n1026 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U721  ( .A0(\U1/aes_core/SB0/n291 ), 
        .A1(\U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n147 ), .B1(
        \U1/aes_core/SB0/n241 ), .C0(\U1/aes_core/SB0/n133 ), .C1(
        \U1/aes_core/SB0/n190 ), .Y(\U1/aes_core/SB0/n1027 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U720  ( .A(\U1/aes_core/SB0/n98 ), .B(
        \U1/aes_core/SB0/n1032 ), .Y(\U1/aes_core/SB0/n327 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U719  ( .A(\U1/aes_core/SB0/n111 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n320 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U718  ( .A(\U1/aes_core/SB0/n169 ), .B(
        \U1/aes_core/SB0/n116 ), .Y(\U1/aes_core/SB0/n310 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U717  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n101 ), .Y(\U1/aes_core/SB0/n206 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U716  ( .AN(\U1/aes_core/SB0/n327 ), .B(
        \U1/aes_core/SB0/n320 ), .C(\U1/aes_core/SB0/n310 ), .D(
        \U1/aes_core/SB0/n206 ), .Y(\U1/aes_core/SB0/n1028 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U715  ( .A(\U1/aes_core/SB0/n209 ), .B(
        \U1/aes_core/SB0/n1031 ), .Y(\U1/aes_core/SB0/n227 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U714  ( .A(\U1/aes_core/SB0/n131 ), .B(
        \U1/aes_core/SB0/n147 ), .Y(\U1/aes_core/SB0/n174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U712  ( .A(\U1/aes_core/SB0/n387 ), .B(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n361 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U710  ( .A(\U1/aes_core/SB0/n386 ), .B(
        \U1/aes_core/SB0/n1025 ), .C(\U1/aes_core/SB0/n1026 ), .D(
        \U1/aes_core/SB0/n1027 ), .E(\U1/aes_core/SB0/n1028 ), .F(
        \U1/aes_core/SB0/n1029 ), .Y(\U1/aes_core/SB0/n451 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U709  ( .A(\U1/aes_core/SB0/n193 ), .B(
        \U1/aes_core/SB0/n371 ), .Y(\U1/aes_core/SB0/n373 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U708  ( .A(\U1/aes_core/SB0/n241 ), .B(
        \U1/aes_core/SB0/n291 ), .Y(\U1/aes_core/SB0/n161 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U707  ( .A(\U1/aes_core/SB0/n260 ), .B(
        \U1/aes_core/SB0/n190 ), .Y(\U1/aes_core/SB0/n323 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U706  ( .A(\U1/aes_core/SB0/n96 ), .B(
        \U1/aes_core/SB0/n190 ), .Y(\U1/aes_core/SB0/n308 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U705  ( .A(\U1/aes_core/SB0/n165 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U704  ( .A(\U1/aes_core/SB0/n115 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n356 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U703  ( .A(\U1/aes_core/SB0/n111 ), .B(
        \U1/aes_core/SB0/n115 ), .Y(\U1/aes_core/SB0/n262 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U702  ( .A(\U1/aes_core/SB0/n201 ), .B(
        \U1/aes_core/SB0/n144 ), .Y(\U1/aes_core/SB0/n337 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U701  ( .A(\U1/aes_core/SB0/n248 ), .B(
        \U1/aes_core/SB0/n356 ), .C(\U1/aes_core/SB0/n262 ), .D(
        \U1/aes_core/SB0/n337 ), .Y(\U1/aes_core/SB0/n1021 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U700  ( .A(\U1/aes_core/SB0/n96 ), .B(
        \U1/aes_core/SB0/n275 ), .Y(\U1/aes_core/SB0/n287 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U699  ( .A(\U1/aes_core/SB0/n97 ), .B(
        \U1/aes_core/SB0/n291 ), .Y(\U1/aes_core/SB0/n187 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U698  ( .A(\U1/aes_core/SB0/n170 ), .B(
        \U1/aes_core/SB0/n131 ), .Y(\U1/aes_core/SB0/n237 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U697  ( .A(\U1/aes_core/SB0/n209 ), .B(
        \U1/aes_core/SB0/n131 ), .Y(\U1/aes_core/SB0/n388 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U696  ( .A0(\U1/aes_core/SB0/n131 ), .A1(
        \U1/aes_core/SB0/n96 ), .B0(\U1/aes_core/SB0/n275 ), .B1(
        \U1/aes_core/SB0/n170 ), .Y(\U1/aes_core/SB0/n1023 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U695  ( .A0(\U1/aes_core/SB0/n291 ), .A1(
        \U1/aes_core/SB0/n99 ), .B0(\U1/aes_core/SB0/n278 ), .B1(
        \U1/aes_core/SB0/n241 ), .Y(\U1/aes_core/SB0/n1024 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U694  ( .A(\U1/aes_core/SB0/n287 ), .B(
        \U1/aes_core/SB0/n187 ), .C(\U1/aes_core/SB0/n237 ), .D(
        \U1/aes_core/SB0/n388 ), .E(\U1/aes_core/SB0/n1023 ), .F(
        \U1/aes_core/SB0/n1024 ), .Y(\U1/aes_core/SB0/n1022 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U693  ( .A(\U1/aes_core/SB0/n373 ), .B(
        \U1/aes_core/SB0/n161 ), .C(\U1/aes_core/SB0/n323 ), .D(
        \U1/aes_core/SB0/n308 ), .E(\U1/aes_core/SB0/n1021 ), .F(
        \U1/aes_core/SB0/n1022 ), .Y(\U1/aes_core/SB0/n462 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U692  ( .A0(\U1/aes_core/SB0/n165 ), 
        .A1(\U1/aes_core/SB0/n168 ), .B0(\U1/aes_core/SB0/n112 ), .B1(
        \U1/aes_core/SB0/n224 ), .C0(\U1/aes_core/SB0/n462 ), .Y(
        \U1/aes_core/SB0/n1020 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U691  ( .A(\U1/aes_core/SB0/n1020 ), .Y(
        \U1/aes_core/SB0/n1013 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U690  ( .A(\U1/aes_core/SB0/n133 ), .B(
        \U1/aes_core/SB0/n170 ), .Y(\U1/aes_core/SB0/n143 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U689  ( .A0(\U1/aes_core/SB0/n166 ), .A1(
        \U1/aes_core/SB0/n143 ), .B0(\U1/aes_core/SB0/n111 ), .Y(
        \U1/aes_core/SB0/n1017 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U688  ( .A0(\U1/aes_core/SB0/n201 ), .A1(
        \U1/aes_core/SB0/n122 ), .B0(\U1/aes_core/SB0/n159 ), .Y(
        \U1/aes_core/SB0/n1018 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U687  ( .A0(\U1/aes_core/SB0/n202 ), .A1(
        \U1/aes_core/SB0/n160 ), .B0(\U1/aes_core/SB0/n116 ), .Y(
        \U1/aes_core/SB0/n1019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U686  ( .A(\U1/aes_core/SB0/n169 ), .B(
        \U1/aes_core/SB0/n123 ), .Y(\U1/aes_core/SB0/n344 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U685  ( .A(\U1/aes_core/SB0/n1017 ), .B(
        \U1/aes_core/SB0/n1018 ), .C(\U1/aes_core/SB0/n1019 ), .D(
        \U1/aes_core/SB0/n344 ), .Y(\U1/aes_core/SB0/n1014 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U684  ( .A(\U1/aes_core/SB0/n124 ), .B(
        \U1/aes_core/SB0/n208 ), .Y(\U1/aes_core/SB0/n154 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB0/U683  ( .A(\U1/aes_core/SB0/n154 ), .B(
        \U1/aes_core/SB0/n134 ), .C(\U1/aes_core/SB0/n147 ), .Y(
        \U1/aes_core/SB0/n1016 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U682  ( .A0(\U1/aes_core/SB0/n170 ), 
        .A1(\U1/aes_core/SB0/n97 ), .B0(\U1/aes_core/SB0/n1016 ), .B1(
        \U1/aes_core/SB0/n136 ), .C0(\U1/aes_core/SB0/n98 ), .C1(
        \U1/aes_core/SB0/n106 ), .Y(\U1/aes_core/SB0/n1015 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U681  ( .A(\U1/aes_core/SB0/n91 ), .B(
        \U1/aes_core/SB0/n451 ), .C(\U1/aes_core/SB0/n1012 ), .D(
        \U1/aes_core/SB0/n1013 ), .E(\U1/aes_core/SB0/n1014 ), .F(
        \U1/aes_core/SB0/n1015 ), .Y(\U1/aes_core/sb0 [1]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U680  ( .A0(\U1/aes_core/SB0/n997 ), .A1(
        \U1/aes_core/SB0/n882 ), .B0(\U1/aes_core/SB0/n938 ), .Y(
        \U1/aes_core/SB0/n1000 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U679  ( .A(\U1/aes_core/SB0/n1009 ), .B(
        \U1/aes_core/SB0/n1010 ), .C(\U1/aes_core/SB0/n1011 ), .Y(
        \U1/aes_core/SB0/n1001 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U678  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n859 ), .Y(\U1/aes_core/SB0/n1006 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U677  ( .A(\U1/aes_core/SB0/n888 ), .B(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n1008 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U676  ( .A0(\U1/aes_core/SB0/n1006 ), 
        .A1(\U1/aes_core/SB0/n1007 ), .B0(\U1/aes_core/SB0/n1008 ), .B1(
        \U1/aes_core/SB0/n865 ), .C0(\U1/aes_core/SB0/n882 ), .C1(
        \U1/aes_core/SB0/n956 ), .Y(\U1/aes_core/SB0/n1002 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U675  ( .A0(\U1/aes_core/SB0/n905 ), 
        .A1(\U1/aes_core/SB0/n1004 ), .B0(\U1/aes_core/SB0/n843 ), .B1(
        \U1/aes_core/SB0/n853 ), .C0(\U1/aes_core/SB0/n880 ), .C1(
        \U1/aes_core/SB0/n1005 ), .Y(\U1/aes_core/SB0/n1003 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U674  ( .A(\U1/aes_core/SB0/n998 ), .B(
        \U1/aes_core/SB0/n999 ), .C(\U1/aes_core/SB0/n1000 ), .D(
        \U1/aes_core/SB0/n1001 ), .E(\U1/aes_core/SB0/n1002 ), .F(
        \U1/aes_core/SB0/n1003 ), .Y(\U1/aes_core/SB0/n873 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U673  ( .A0(\U1/aes_core/SB0/n997 ), .A1(
        \U1/aes_core/SB0/n988 ), .B0(\U1/aes_core/SB0/n917 ), .Y(
        \U1/aes_core/SB0/n962 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB0/U672  ( .A0(\U1/aes_core/SB0/n893 ), .A1(
        \U1/aes_core/SB0/n880 ), .A2(\U1/aes_core/SB0/n940 ), .B0(
        \U1/aes_core/SB0/n864 ), .Y(\U1/aes_core/SB0/n963 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U671  ( .A(\U1/aes_core/SB0/n993 ), .B(
        \U1/aes_core/SB0/n994 ), .C(\U1/aes_core/SB0/n995 ), .D(
        \U1/aes_core/SB0/n996 ), .Y(\U1/aes_core/SB0/n966 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U670  ( .A(\U1/aes_core/SB0/n992 ), .Y(
        \U1/aes_core/SB0/n969 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U669  ( .A(\U1/aes_core/SB0/n991 ), .Y(
        \U1/aes_core/SB0/n975 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB0/U668  ( .A0(\U1/aes_core/SB0/n989 ), 
        .A1(\U1/aes_core/SB0/n852 ), .B0N(\U1/aes_core/SB0/n990 ), .Y(
        \U1/aes_core/SB0/n976 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U667  ( .A0(\U1/aes_core/SB0/n845 ), 
        .A1(\U1/aes_core/SB0/n988 ), .B0(\U1/aes_core/SB0/n938 ), .B1(
        \U1/aes_core/SB0/n878 ), .C0(\U1/aes_core/SB0/n864 ), .C1(
        \U1/aes_core/SB0/n843 ), .Y(\U1/aes_core/SB0/n977 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U666  ( .AN(\U1/aes_core/SB0/n984 ), .B(
        \U1/aes_core/SB0/n985 ), .C(\U1/aes_core/SB0/n986 ), .D(
        \U1/aes_core/SB0/n987 ), .Y(\U1/aes_core/SB0/n978 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U665  ( .A(\U1/aes_core/SB0/n980 ), .B(
        \U1/aes_core/SB0/n981 ), .C(\U1/aes_core/SB0/n982 ), .D(
        \U1/aes_core/SB0/n983 ), .Y(\U1/aes_core/SB0/n979 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U664  ( .A(\U1/aes_core/SB0/n974 ), .B(
        \U1/aes_core/SB0/n975 ), .C(\U1/aes_core/SB0/n976 ), .D(
        \U1/aes_core/SB0/n977 ), .E(\U1/aes_core/SB0/n978 ), .F(
        \U1/aes_core/SB0/n979 ), .Y(\U1/aes_core/SB0/n973 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U663  ( .A(\U1/aes_core/SB0/n973 ), .Y(
        \U1/aes_core/SB0/n895 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U662  ( .A0(\U1/aes_core/SB0/n905 ), .A1(
        \U1/aes_core/SB0/n883 ), .B0(\U1/aes_core/SB0/n843 ), .B1(
        \U1/aes_core/SB0/n844 ), .Y(\U1/aes_core/SB0/n972 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U661  ( .A0(\U1/aes_core/SB0/n915 ), 
        .A1(\U1/aes_core/SB0/n971 ), .B0(\U1/aes_core/SB0/n891 ), .B1(
        \U1/aes_core/SB0/n869 ), .C0(\U1/aes_core/SB0/n972 ), .Y(
        \U1/aes_core/SB0/n970 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U660  ( .AN(\U1/aes_core/SB0/n968 ), .B(
        \U1/aes_core/SB0/n969 ), .C(\U1/aes_core/SB0/n895 ), .D(
        \U1/aes_core/SB0/n970 ), .Y(\U1/aes_core/SB0/n967 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U659  ( .A(\U1/aes_core/SB0/n962 ), .B(
        \U1/aes_core/SB0/n963 ), .C(\U1/aes_core/SB0/n964 ), .D(
        \U1/aes_core/SB0/n965 ), .E(\U1/aes_core/SB0/n966 ), .F(
        \U1/aes_core/SB0/n967 ), .Y(\U1/aes_core/SB0/n897 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U658  ( .A(\U1/aes_core/SB0/n961 ), .Y(
        \U1/aes_core/SB0/n957 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U657  ( .A0(\U1/aes_core/SB0/n959 ), .A1(
        \U1/aes_core/SB0/n960 ), .B0(\U1/aes_core/SB0/n913 ), .B1(
        \U1/aes_core/SB0/n954 ), .Y(\U1/aes_core/SB0/n958 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U656  ( .A0(\U1/aes_core/SB0/n864 ), 
        .A1(\U1/aes_core/SB0/n956 ), .B0(\U1/aes_core/SB0/n957 ), .C0(
        \U1/aes_core/SB0/n958 ), .Y(\U1/aes_core/SB0/n942 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U655  ( .A0(\U1/aes_core/SB0/n955 ), .A1(
        \U1/aes_core/SB0/n892 ), .B0(\U1/aes_core/SB0/n863 ), .Y(
        \U1/aes_core/SB0/n950 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U654  ( .A0(\U1/aes_core/SB0/n954 ), .A1(
        \U1/aes_core/SB0/n889 ), .B0(\U1/aes_core/SB0/n860 ), .Y(
        \U1/aes_core/SB0/n951 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U653  ( .A(\U1/aes_core/SB0/n950 ), .B(
        \U1/aes_core/SB0/n951 ), .C(\U1/aes_core/SB0/n952 ), .D(
        \U1/aes_core/SB0/n953 ), .Y(\U1/aes_core/SB0/n943 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U652  ( .A(\U1/aes_core/SB0/n912 ), .B(
        \U1/aes_core/SB0/n949 ), .Y(\U1/aes_core/SB0/n945 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U651  ( .A(\U1/aes_core/SB0/n948 ), .B(
        \U1/aes_core/SB0/n907 ), .Y(\U1/aes_core/SB0/n946 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U650  ( .A0(\U1/aes_core/SB0/n945 ), 
        .A1(\U1/aes_core/SB0/n846 ), .B0(\U1/aes_core/SB0/n946 ), .B1(
        \U1/aes_core/SB0/n882 ), .C0(\U1/aes_core/SB0/n947 ), .C1(
        \U1/aes_core/SB0/n881 ), .Y(\U1/aes_core/SB0/n944 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U649  ( .A(\U1/aes_core/SB0/n873 ), .B(
        \U1/aes_core/SB0/n897 ), .C(\U1/aes_core/SB0/n941 ), .D(
        \U1/aes_core/SB0/n942 ), .E(\U1/aes_core/SB0/n943 ), .F(
        \U1/aes_core/SB0/n944 ), .Y(\U1/aes_core/sb0 [20]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U648  ( .A1N(\U1/aes_core/SB0/n939 ), 
        .A0(\U1/aes_core/SB0/n940 ), .B0(\U1/aes_core/SB0/n883 ), .Y(
        \U1/aes_core/SB0/n923 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U647  ( .A(\U1/aes_core/SB0/n870 ), .B(
        \U1/aes_core/SB0/n889 ), .Y(\U1/aes_core/SB0/n936 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U646  ( .A0(\U1/aes_core/SB0/n846 ), 
        .A1(\U1/aes_core/SB0/n935 ), .B0(\U1/aes_core/SB0/n936 ), .B1(
        \U1/aes_core/SB0/n843 ), .C0(\U1/aes_core/SB0/n937 ), .C1(
        \U1/aes_core/SB0/n938 ), .Y(\U1/aes_core/SB0/n924 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U645  ( .A(\U1/aes_core/SB0/n934 ), .Y(
        \U1/aes_core/SB0/n931 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U644  ( .AN(\U1/aes_core/SB0/n930 ), .B(
        \U1/aes_core/SB0/n931 ), .C(\U1/aes_core/SB0/n932 ), .D(
        \U1/aes_core/SB0/n933 ), .Y(\U1/aes_core/SB0/n925 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U643  ( .A(\U1/aes_core/SB0/n927 ), .B(
        \U1/aes_core/SB0/n928 ), .C(\U1/aes_core/SB0/n929 ), .Y(
        \U1/aes_core/SB0/n926 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U642  ( .A(\U1/aes_core/SB0/n921 ), .B(
        \U1/aes_core/SB0/n922 ), .C(\U1/aes_core/SB0/n923 ), .D(
        \U1/aes_core/SB0/n924 ), .E(\U1/aes_core/SB0/n925 ), .F(
        \U1/aes_core/SB0/n926 ), .Y(\U1/aes_core/SB0/n872 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U641  ( .A(\U1/aes_core/SB0/n920 ), .Y(
        \U1/aes_core/SB0/n918 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U640  ( .A0(\U1/aes_core/SB0/n859 ), .A1(
        \U1/aes_core/SB0/n862 ), .B0(\U1/aes_core/SB0/n858 ), .B1(
        \U1/aes_core/SB0/n860 ), .Y(\U1/aes_core/SB0/n919 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U639  ( .A0(\U1/aes_core/SB0/n883 ), 
        .A1(\U1/aes_core/SB0/n917 ), .B0(\U1/aes_core/SB0/n918 ), .C0(
        \U1/aes_core/SB0/n919 ), .Y(\U1/aes_core/SB0/n898 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U638  ( .A0(\U1/aes_core/SB0/n915 ), .A1(
        \U1/aes_core/SB0/n859 ), .B0(\U1/aes_core/SB0/n916 ), .Y(
        \U1/aes_core/SB0/n909 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U637  ( .A0(\U1/aes_core/SB0/n912 ), .A1(
        \U1/aes_core/SB0/n913 ), .B0(\U1/aes_core/SB0/n914 ), .Y(
        \U1/aes_core/SB0/n910 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U636  ( .AN(\U1/aes_core/SB0/n908 ), .B(
        \U1/aes_core/SB0/n909 ), .C(\U1/aes_core/SB0/n910 ), .D(
        \U1/aes_core/SB0/n911 ), .Y(\U1/aes_core/SB0/n899 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U635  ( .A0(\U1/aes_core/SB0/n863 ), .A1(
        \U1/aes_core/SB0/n906 ), .B0(\U1/aes_core/SB0/n907 ), .Y(
        \U1/aes_core/SB0/n902 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB0/U634  ( .A0(\U1/aes_core/SB0/n881 ), .A1(
        \U1/aes_core/SB0/n904 ), .B0(\U1/aes_core/SB0/n844 ), .B1(
        \U1/aes_core/SB0/n905 ), .Y(\U1/aes_core/SB0/n903 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U633  ( .A0(\U1/aes_core/SB0/n901 ), 
        .A1(\U1/aes_core/SB0/n882 ), .B0(\U1/aes_core/SB0/n902 ), .C0(
        \U1/aes_core/SB0/n903 ), .Y(\U1/aes_core/SB0/n900 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U632  ( .A(\U1/aes_core/SB0/n872 ), .B(
        \U1/aes_core/SB0/n896 ), .C(\U1/aes_core/SB0/n897 ), .D(
        \U1/aes_core/SB0/n898 ), .E(\U1/aes_core/SB0/n899 ), .F(
        \U1/aes_core/SB0/n900 ), .Y(\U1/aes_core/sb0 [21]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U631  ( .A0(\U1/aes_core/SB0/n893 ), 
        .A1(\U1/aes_core/SB0/n853 ), .B0(\U1/aes_core/SB0/n894 ), .B1(
        \U1/aes_core/SB0/n846 ), .C0(\U1/aes_core/SB0/n895 ), .Y(
        \U1/aes_core/SB0/n875 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U630  ( .A0(\U1/aes_core/SB0/n892 ), .A1(
        \U1/aes_core/SB0/n848 ), .B0(\U1/aes_core/SB0/n859 ), .Y(
        \U1/aes_core/SB0/n884 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U629  ( .A0(\U1/aes_core/SB0/n868 ), .A1(
        \U1/aes_core/SB0/n891 ), .B0(\U1/aes_core/SB0/n860 ), .Y(
        \U1/aes_core/SB0/n885 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U628  ( .A0(\U1/aes_core/SB0/n888 ), .A1(
        \U1/aes_core/SB0/n889 ), .B0(\U1/aes_core/SB0/n890 ), .Y(
        \U1/aes_core/SB0/n886 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U627  ( .A(\U1/aes_core/SB0/n884 ), .B(
        \U1/aes_core/SB0/n885 ), .C(\U1/aes_core/SB0/n886 ), .D(
        \U1/aes_core/SB0/n887 ), .Y(\U1/aes_core/SB0/n876 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U626  ( .A(\U1/aes_core/SB0/n853 ), .B(
        \U1/aes_core/SB0/n883 ), .Y(\U1/aes_core/SB0/n851 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U625  ( .A(\U1/aes_core/SB0/n863 ), .B(
        \U1/aes_core/SB0/n851 ), .Y(\U1/aes_core/SB0/n879 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U624  ( .A0(\U1/aes_core/SB0/n865 ), 
        .A1(\U1/aes_core/SB0/n878 ), .B0(\U1/aes_core/SB0/n879 ), .B1(
        \U1/aes_core/SB0/n880 ), .C0(\U1/aes_core/SB0/n881 ), .C1(
        \U1/aes_core/SB0/n882 ), .Y(\U1/aes_core/SB0/n877 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U623  ( .A(\U1/aes_core/SB0/n872 ), .B(
        \U1/aes_core/SB0/n873 ), .C(\U1/aes_core/SB0/n874 ), .D(
        \U1/aes_core/SB0/n875 ), .E(\U1/aes_core/SB0/n876 ), .F(
        \U1/aes_core/SB0/n877 ), .Y(\U1/aes_core/sb0 [22]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U622  ( .A0(\U1/aes_core/SB0/n868 ), .A1(
        \U1/aes_core/SB0/n869 ), .B0(\U1/aes_core/SB0/n870 ), .B1(
        \U1/aes_core/SB0/n871 ), .Y(\U1/aes_core/SB0/n867 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U621  ( .A0(\U1/aes_core/SB0/n864 ), 
        .A1(\U1/aes_core/SB0/n865 ), .B0(\U1/aes_core/SB0/n866 ), .C0(
        \U1/aes_core/SB0/n867 ), .Y(\U1/aes_core/SB0/n840 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U620  ( .A1N(\U1/aes_core/SB0/n861 ), 
        .A0(\U1/aes_core/SB0/n862 ), .B0(\U1/aes_core/SB0/n863 ), .Y(
        \U1/aes_core/SB0/n854 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U619  ( .A0(\U1/aes_core/SB0/n858 ), .A1(
        \U1/aes_core/SB0/n859 ), .B0(\U1/aes_core/SB0/n860 ), .Y(
        \U1/aes_core/SB0/n855 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U618  ( .A(\U1/aes_core/SB0/n854 ), .B(
        \U1/aes_core/SB0/n855 ), .C(\U1/aes_core/SB0/n856 ), .D(
        \U1/aes_core/SB0/n857 ), .Y(\U1/aes_core/SB0/n841 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U617  ( .A(\U1/aes_core/SB0/n852 ), .B(
        \U1/aes_core/SB0/n853 ), .Y(\U1/aes_core/SB0/n849 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U616  ( .A0(\U1/aes_core/SB0/n848 ), .A1(
        \U1/aes_core/SB0/n849 ), .B0(\U1/aes_core/SB0/n850 ), .B1(
        \U1/aes_core/SB0/n851 ), .Y(\U1/aes_core/SB0/n847 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U615  ( .A0(\U1/aes_core/SB0/n843 ), 
        .A1(\U1/aes_core/SB0/n844 ), .B0(\U1/aes_core/SB0/n845 ), .B1(
        \U1/aes_core/SB0/n846 ), .C0(\U1/aes_core/SB0/n847 ), .Y(
        \U1/aes_core/SB0/n842 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U614  ( .A(\U1/aes_core/SB0/n837 ), .B(
        \U1/aes_core/SB0/n838 ), .C(\U1/aes_core/SB0/n839 ), .D(
        \U1/aes_core/SB0/n840 ), .E(\U1/aes_core/SB0/n841 ), .F(
        \U1/aes_core/SB0/n842 ), .Y(\U1/aes_core/sb0 [23]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U613  ( .A(Dout[127]), .B(Dout[126]), .Y(
        \U1/aes_core/SB0/n818 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U612  ( .A(Dout[125]), .B(Dout[124]), .Y(
        \U1/aes_core/SB0/n827 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U611  ( .A(\U1/aes_core/SB0/n818 ), .B(
        \U1/aes_core/SB0/n827 ), .Y(\U1/aes_core/SB0/n753 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U610  ( .A(Dout[121]), .Y(
        \U1/aes_core/SB0/n833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U609  ( .A(Dout[120]), .Y(
        \U1/aes_core/SB0/n836 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U608  ( .A(\U1/aes_core/SB0/n833 ), .B(
        \U1/aes_core/SB0/n836 ), .Y(\U1/aes_core/SB0/n826 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U607  ( .A(Dout[123]), .B(Dout[122]), .Y(
        \U1/aes_core/SB0/n806 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U606  ( .A(\U1/aes_core/SB0/n826 ), .B(
        \U1/aes_core/SB0/n806 ), .Y(\U1/aes_core/SB0/n448 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U605  ( .A(\U1/aes_core/SB0/n753 ), .B(
        \U1/aes_core/SB0/n448 ), .Y(\U1/aes_core/SB0/n662 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U604  ( .A(Dout[122]), .B(Dout[123]), .Y(
        \U1/aes_core/SB0/n823 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U603  ( .A(\U1/aes_core/SB0/n823 ), .B(
        \U1/aes_core/SB0/n826 ), .Y(\U1/aes_core/SB0/n531 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U602  ( .A(Dout[127]), .Y(
        \U1/aes_core/SB0/n830 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U601  ( .A(\U1/aes_core/SB0/n830 ), .B(
        Dout[126]), .Y(\U1/aes_core/SB0/n800 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U600  ( .A(\U1/aes_core/SB0/n800 ), .B(
        \U1/aes_core/SB0/n827 ), .Y(\U1/aes_core/SB0/n754 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U599  ( .A(\U1/aes_core/SB0/n531 ), .B(
        \U1/aes_core/SB0/n754 ), .Y(\U1/aes_core/SB0/n565 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U598  ( .A(Dout[123]), .Y(
        \U1/aes_core/SB0/n835 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB0/U597  ( .A(Dout[122]), .B(
        \U1/aes_core/SB0/n835 ), .Y(\U1/aes_core/SB0/n825 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U596  ( .A(\U1/aes_core/SB0/n826 ), .B(
        \U1/aes_core/SB0/n825 ), .Y(\U1/aes_core/SB0/n600 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U595  ( .A(\U1/aes_core/SB0/n600 ), .Y(
        \U1/aes_core/SB0/n414 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U594  ( .A(Dout[124]), .Y(
        \U1/aes_core/SB0/n834 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U593  ( .A(\U1/aes_core/SB0/n834 ), .B(
        Dout[125]), .Y(\U1/aes_core/SB0/n819 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U592  ( .A(Dout[126]), .Y(
        \U1/aes_core/SB0/n831 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U591  ( .A(\U1/aes_core/SB0/n831 ), .B(
        Dout[127]), .Y(\U1/aes_core/SB0/n809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U590  ( .A(\U1/aes_core/SB0/n819 ), .B(
        \U1/aes_core/SB0/n809 ), .Y(\U1/aes_core/SB0/n579 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U589  ( .A(\U1/aes_core/SB0/n579 ), .Y(
        \U1/aes_core/SB0/n481 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U588  ( .A(\U1/aes_core/SB0/n414 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n622 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U587  ( .A(\U1/aes_core/SB0/n753 ), .Y(
        \U1/aes_core/SB0/n445 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U586  ( .A(Dout[121]), .B(Dout[120]), .Y(
        \U1/aes_core/SB0/n822 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U585  ( .A(\U1/aes_core/SB0/n822 ), .B(
        \U1/aes_core/SB0/n806 ), .Y(\U1/aes_core/SB0/n513 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U584  ( .A(\U1/aes_core/SB0/n513 ), .Y(
        \U1/aes_core/SB0/n404 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U583  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n404 ), .Y(\U1/aes_core/SB0/n508 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U582  ( .A(\U1/aes_core/SB0/n836 ), .B(
        Dout[121]), .Y(\U1/aes_core/SB0/n807 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U581  ( .A(\U1/aes_core/SB0/n825 ), .B(
        \U1/aes_core/SB0/n807 ), .Y(\U1/aes_core/SB0/n613 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U580  ( .A(\U1/aes_core/SB0/n613 ), .Y(
        \U1/aes_core/SB0/n524 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U579  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n644 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U578  ( .A(\U1/aes_core/SB0/n622 ), .B(
        \U1/aes_core/SB0/n508 ), .C(\U1/aes_core/SB0/n644 ), .Y(
        \U1/aes_core/SB0/n787 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U577  ( .A(\U1/aes_core/SB0/n827 ), .B(
        \U1/aes_core/SB0/n809 ), .Y(\U1/aes_core/SB0/n580 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U576  ( .A(\U1/aes_core/SB0/n835 ), .B(
        Dout[122]), .Y(\U1/aes_core/SB0/n816 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U575  ( .A(\U1/aes_core/SB0/n816 ), .B(
        \U1/aes_core/SB0/n807 ), .Y(\U1/aes_core/SB0/n582 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U574  ( .A(\U1/aes_core/SB0/n580 ), .B(
        \U1/aes_core/SB0/n582 ), .Y(\U1/aes_core/SB0/n667 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U573  ( .A(\U1/aes_core/SB0/n754 ), .Y(
        \U1/aes_core/SB0/n443 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U572  ( .A(Dout[125]), .Y(
        \U1/aes_core/SB0/n832 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U571  ( .A(\U1/aes_core/SB0/n834 ), .B(
        \U1/aes_core/SB0/n832 ), .Y(\U1/aes_core/SB0/n808 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U570  ( .A(\U1/aes_core/SB0/n818 ), .B(
        \U1/aes_core/SB0/n808 ), .Y(\U1/aes_core/SB0/n400 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U569  ( .A(\U1/aes_core/SB0/n400 ), .Y(
        \U1/aes_core/SB0/n490 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U568  ( .A(\U1/aes_core/SB0/n833 ), .B(
        Dout[120]), .Y(\U1/aes_core/SB0/n817 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U567  ( .A(\U1/aes_core/SB0/n817 ), .B(
        \U1/aes_core/SB0/n806 ), .Y(\U1/aes_core/SB0/n435 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U566  ( .A(\U1/aes_core/SB0/n435 ), .Y(
        \U1/aes_core/SB0/n608 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U565  ( .A0(\U1/aes_core/SB0/n443 ), .A1(
        \U1/aes_core/SB0/n490 ), .B0(\U1/aes_core/SB0/n608 ), .Y(
        \U1/aes_core/SB0/n828 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U564  ( .A(\U1/aes_core/SB0/n822 ), .B(
        \U1/aes_core/SB0/n825 ), .Y(\U1/aes_core/SB0/n447 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U563  ( .A(\U1/aes_core/SB0/n447 ), .Y(
        \U1/aes_core/SB0/n482 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U562  ( .A(\U1/aes_core/SB0/n832 ), .B(
        Dout[124]), .Y(\U1/aes_core/SB0/n801 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U561  ( .A(\U1/aes_core/SB0/n809 ), .B(
        \U1/aes_core/SB0/n801 ), .Y(\U1/aes_core/SB0/n407 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U560  ( .A(\U1/aes_core/SB0/n580 ), .B(
        \U1/aes_core/SB0/n407 ), .Y(\U1/aes_core/SB0/n689 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U559  ( .A(\U1/aes_core/SB0/n830 ), .B(
        \U1/aes_core/SB0/n831 ), .Y(\U1/aes_core/SB0/n810 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U558  ( .A(\U1/aes_core/SB0/n819 ), .B(
        \U1/aes_core/SB0/n810 ), .Y(\U1/aes_core/SB0/n432 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U557  ( .A(\U1/aes_core/SB0/n432 ), .Y(
        \U1/aes_core/SB0/n709 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U556  ( .A0(\U1/aes_core/SB0/n482 ), .A1(
        \U1/aes_core/SB0/n689 ), .B0(\U1/aes_core/SB0/n709 ), .B1(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n829 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U555  ( .AN(\U1/aes_core/SB0/n667 ), .B(
        \U1/aes_core/SB0/n828 ), .C(\U1/aes_core/SB0/n829 ), .Y(
        \U1/aes_core/SB0/n788 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U554  ( .A(\U1/aes_core/SB0/n827 ), .B(
        \U1/aes_core/SB0/n810 ), .Y(\U1/aes_core/SB0/n563 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U553  ( .A(\U1/aes_core/SB0/n823 ), .B(
        \U1/aes_core/SB0/n822 ), .Y(\U1/aes_core/SB0/n397 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U552  ( .A(\U1/aes_core/SB0/n800 ), .B(
        \U1/aes_core/SB0/n819 ), .Y(\U1/aes_core/SB0/n512 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U551  ( .A(\U1/aes_core/SB0/n823 ), .B(
        \U1/aes_core/SB0/n817 ), .Y(\U1/aes_core/SB0/n515 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U550  ( .A(\U1/aes_core/SB0/n826 ), .B(
        \U1/aes_core/SB0/n816 ), .Y(\U1/aes_core/SB0/n510 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U549  ( .A(\U1/aes_core/SB0/n510 ), .Y(
        \U1/aes_core/SB0/n530 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U548  ( .A(\U1/aes_core/SB0/n407 ), .Y(
        \U1/aes_core/SB0/n694 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U547  ( .A(\U1/aes_core/SB0/n825 ), .B(
        \U1/aes_core/SB0/n817 ), .Y(\U1/aes_core/SB0/n492 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U546  ( .A(\U1/aes_core/SB0/n492 ), .Y(
        \U1/aes_core/SB0/n446 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U545  ( .A0(\U1/aes_core/SB0/n530 ), .A1(
        \U1/aes_core/SB0/n445 ), .B0(\U1/aes_core/SB0/n694 ), .B1(
        \U1/aes_core/SB0/n446 ), .Y(\U1/aes_core/SB0/n824 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U544  ( .A0(\U1/aes_core/SB0/n563 ), 
        .A1(\U1/aes_core/SB0/n397 ), .B0(\U1/aes_core/SB0/n512 ), .B1(
        \U1/aes_core/SB0/n515 ), .C0(\U1/aes_core/SB0/n824 ), .Y(
        \U1/aes_core/SB0/n789 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U543  ( .A(\U1/aes_core/SB0/n510 ), .B(
        \U1/aes_core/SB0/n563 ), .Y(\U1/aes_core/SB0/n701 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U542  ( .A(\U1/aes_core/SB0/n515 ), .B(
        \U1/aes_core/SB0/n580 ), .Y(\U1/aes_core/SB0/n691 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U541  ( .A(\U1/aes_core/SB0/n691 ), .Y(
        \U1/aes_core/SB0/n820 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U540  ( .A(\U1/aes_core/SB0/n823 ), .B(
        \U1/aes_core/SB0/n807 ), .Y(\U1/aes_core/SB0/n419 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U539  ( .A(\U1/aes_core/SB0/n419 ), .Y(
        \U1/aes_core/SB0/n491 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U538  ( .A(\U1/aes_core/SB0/n822 ), .B(
        \U1/aes_core/SB0/n816 ), .Y(\U1/aes_core/SB0/n434 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U537  ( .A(\U1/aes_core/SB0/n434 ), .Y(
        \U1/aes_core/SB0/n423 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U536  ( .A0(\U1/aes_core/SB0/n491 ), .A1(
        \U1/aes_core/SB0/n423 ), .B0(\U1/aes_core/SB0/n490 ), .Y(
        \U1/aes_core/SB0/n821 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U535  ( .A(\U1/aes_core/SB0/n818 ), .B(
        \U1/aes_core/SB0/n801 ), .Y(\U1/aes_core/SB0/n418 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U534  ( .A(\U1/aes_core/SB0/n418 ), .Y(
        \U1/aes_core/SB0/n489 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U533  ( .A(\U1/aes_core/SB0/n489 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n674 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U532  ( .AN(\U1/aes_core/SB0/n701 ), .B(
        \U1/aes_core/SB0/n820 ), .C(\U1/aes_core/SB0/n821 ), .D(
        \U1/aes_core/SB0/n674 ), .Y(\U1/aes_core/SB0/n811 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U531  ( .A(\U1/aes_core/SB0/n808 ), .B(
        \U1/aes_core/SB0/n810 ), .Y(\U1/aes_core/SB0/n398 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U530  ( .A(\U1/aes_core/SB0/n818 ), .B(
        \U1/aes_core/SB0/n819 ), .Y(\U1/aes_core/SB0/n406 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U529  ( .A0(\U1/aes_core/SB0/n754 ), 
        .A1(\U1/aes_core/SB0/n600 ), .B0(\U1/aes_core/SB0/n398 ), .B1(
        \U1/aes_core/SB0/n510 ), .C0(\U1/aes_core/SB0/n406 ), .C1(
        \U1/aes_core/SB0/n492 ), .Y(\U1/aes_core/SB0/n812 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U528  ( .A(\U1/aes_core/SB0/n447 ), .B(
        \U1/aes_core/SB0/n754 ), .Y(\U1/aes_core/SB0/n616 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U527  ( .A(\U1/aes_core/SB0/n694 ), .B(
        \U1/aes_core/SB0/n530 ), .Y(\U1/aes_core/SB0/n663 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U526  ( .A(\U1/aes_core/SB0/n446 ), .B(
        \U1/aes_core/SB0/n445 ), .Y(\U1/aes_core/SB0/n643 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U525  ( .A(\U1/aes_core/SB0/n512 ), .Y(
        \U1/aes_core/SB0/n417 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U524  ( .A(\U1/aes_core/SB0/n417 ), .B(
        \U1/aes_core/SB0/n608 ), .Y(\U1/aes_core/SB0/n605 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U523  ( .AN(\U1/aes_core/SB0/n616 ), .B(
        \U1/aes_core/SB0/n663 ), .C(\U1/aes_core/SB0/n643 ), .D(
        \U1/aes_core/SB0/n605 ), .Y(\U1/aes_core/SB0/n813 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U522  ( .A(\U1/aes_core/SB0/n800 ), .B(
        \U1/aes_core/SB0/n808 ), .Y(\U1/aes_core/SB0/n693 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U521  ( .A(\U1/aes_core/SB0/n693 ), .B(
        \U1/aes_core/SB0/n435 ), .Y(\U1/aes_core/SB0/n539 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U520  ( .A(\U1/aes_core/SB0/n816 ), .B(
        \U1/aes_core/SB0/n817 ), .Y(\U1/aes_core/SB0/n399 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U519  ( .A(\U1/aes_core/SB0/n432 ), .B(
        \U1/aes_core/SB0/n399 ), .Y(\U1/aes_core/SB0/n574 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U518  ( .A(\U1/aes_core/SB0/n574 ), .Y(
        \U1/aes_core/SB0/n815 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U517  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n608 ), .Y(\U1/aes_core/SB0/n555 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U516  ( .A(\U1/aes_core/SB0/n399 ), .Y(
        \U1/aes_core/SB0/n416 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U515  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n416 ), .Y(\U1/aes_core/SB0/n504 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U514  ( .AN(\U1/aes_core/SB0/n539 ), .B(
        \U1/aes_core/SB0/n815 ), .C(\U1/aes_core/SB0/n555 ), .D(
        \U1/aes_core/SB0/n504 ), .Y(\U1/aes_core/SB0/n814 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U513  ( .A(\U1/aes_core/SB0/n811 ), .B(
        \U1/aes_core/SB0/n812 ), .C(\U1/aes_core/SB0/n813 ), .D(
        \U1/aes_core/SB0/n814 ), .Y(\U1/aes_core/SB0/n713 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U512  ( .A(\U1/aes_core/SB0/n513 ), .B(
        \U1/aes_core/SB0/n693 ), .Y(\U1/aes_core/SB0/n505 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U511  ( .A(\U1/aes_core/SB0/n801 ), .B(
        \U1/aes_core/SB0/n810 ), .Y(\U1/aes_core/SB0/n597 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U510  ( .A(\U1/aes_core/SB0/n531 ), .B(
        \U1/aes_core/SB0/n597 ), .Y(\U1/aes_core/SB0/n626 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U509  ( .A(\U1/aes_core/SB0/n398 ), .Y(
        \U1/aes_core/SB0/n442 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U508  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n482 ), .Y(\U1/aes_core/SB0/n677 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U507  ( .A0(\U1/aes_core/SB0/n597 ), .A1(
        \U1/aes_core/SB0/n399 ), .B0(\U1/aes_core/SB0/n677 ), .Y(
        \U1/aes_core/SB0/n802 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U506  ( .A(\U1/aes_core/SB0/n582 ), .Y(
        \U1/aes_core/SB0/n487 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U505  ( .A(\U1/aes_core/SB0/n487 ), .B(
        \U1/aes_core/SB0/n443 ), .Y(\U1/aes_core/SB0/n486 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U504  ( .A(\U1/aes_core/SB0/n443 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n527 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U503  ( .A(\U1/aes_core/SB0/n808 ), .B(
        \U1/aes_core/SB0/n809 ), .Y(\U1/aes_core/SB0/n436 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U502  ( .A(\U1/aes_core/SB0/n436 ), .Y(
        \U1/aes_core/SB0/n682 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U501  ( .A(\U1/aes_core/SB0/n491 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n658 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U500  ( .A(\U1/aes_core/SB0/n448 ), .Y(
        \U1/aes_core/SB0/n488 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U499  ( .A(\U1/aes_core/SB0/n488 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n594 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U498  ( .A(\U1/aes_core/SB0/n486 ), .B(
        \U1/aes_core/SB0/n527 ), .C(\U1/aes_core/SB0/n658 ), .D(
        \U1/aes_core/SB0/n594 ), .Y(\U1/aes_core/SB0/n803 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U497  ( .A(\U1/aes_core/SB0/n446 ), .B(
        \U1/aes_core/SB0/n489 ), .Y(\U1/aes_core/SB0/n560 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U496  ( .A(\U1/aes_core/SB0/n404 ), .B(
        \U1/aes_core/SB0/n489 ), .Y(\U1/aes_core/SB0/n569 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U495  ( .A(\U1/aes_core/SB0/n406 ), .Y(
        \U1/aes_core/SB0/n413 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U494  ( .A(\U1/aes_core/SB0/n530 ), .B(
        \U1/aes_core/SB0/n413 ), .Y(\U1/aes_core/SB0/n697 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U493  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n491 ), .Y(\U1/aes_core/SB0/n586 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U492  ( .A(\U1/aes_core/SB0/n560 ), .B(
        \U1/aes_core/SB0/n569 ), .C(\U1/aes_core/SB0/n697 ), .D(
        \U1/aes_core/SB0/n586 ), .Y(\U1/aes_core/SB0/n804 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U491  ( .A(\U1/aes_core/SB0/n515 ), .Y(
        \U1/aes_core/SB0/n546 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U490  ( .A(\U1/aes_core/SB0/n694 ), .B(
        \U1/aes_core/SB0/n546 ), .Y(\U1/aes_core/SB0/n711 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U489  ( .A(\U1/aes_core/SB0/n806 ), .B(
        \U1/aes_core/SB0/n807 ), .Y(\U1/aes_core/SB0/n480 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U488  ( .A(\U1/aes_core/SB0/n480 ), .Y(
        \U1/aes_core/SB0/n425 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U487  ( .A(\U1/aes_core/SB0/n694 ), .B(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n646 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U486  ( .A(\U1/aes_core/SB0/n531 ), .Y(
        \U1/aes_core/SB0/n402 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U485  ( .A(\U1/aes_core/SB0/n402 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n611 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U484  ( .A(\U1/aes_core/SB0/n490 ), .B(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n441 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U483  ( .A(\U1/aes_core/SB0/n711 ), .B(
        \U1/aes_core/SB0/n646 ), .C(\U1/aes_core/SB0/n611 ), .D(
        \U1/aes_core/SB0/n441 ), .Y(\U1/aes_core/SB0/n805 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U482  ( .A(\U1/aes_core/SB0/n505 ), .B(
        \U1/aes_core/SB0/n626 ), .C(\U1/aes_core/SB0/n802 ), .D(
        \U1/aes_core/SB0/n803 ), .E(\U1/aes_core/SB0/n804 ), .F(
        \U1/aes_core/SB0/n805 ), .Y(\U1/aes_core/SB0/n724 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U481  ( .A(\U1/aes_core/SB0/n724 ), .Y(
        \U1/aes_core/SB0/n791 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U480  ( .A(\U1/aes_core/SB0/n434 ), .B(
        \U1/aes_core/SB0/n597 ), .Y(\U1/aes_core/SB0/n700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U479  ( .A(\U1/aes_core/SB0/n800 ), .B(
        \U1/aes_core/SB0/n801 ), .Y(\U1/aes_core/SB0/n437 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U478  ( .A(\U1/aes_core/SB0/n437 ), .B(
        \U1/aes_core/SB0/n582 ), .Y(\U1/aes_core/SB0/n573 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U477  ( .A(\U1/aes_core/SB0/n573 ), .Y(
        \U1/aes_core/SB0/n798 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U476  ( .A(\U1/aes_core/SB0/n580 ), .Y(
        \U1/aes_core/SB0/n412 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U475  ( .A0(\U1/aes_core/SB0/n682 ), .A1(
        \U1/aes_core/SB0/n412 ), .B0(\U1/aes_core/SB0/n425 ), .Y(
        \U1/aes_core/SB0/n799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U474  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n546 ), .Y(\U1/aes_core/SB0/n675 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U473  ( .AN(\U1/aes_core/SB0/n700 ), .B(
        \U1/aes_core/SB0/n798 ), .C(\U1/aes_core/SB0/n799 ), .D(
        \U1/aes_core/SB0/n675 ), .Y(\U1/aes_core/SB0/n794 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U472  ( .A0(\U1/aes_core/SB0/n448 ), 
        .A1(\U1/aes_core/SB0/n400 ), .B0(\U1/aes_core/SB0/n563 ), .B1(
        \U1/aes_core/SB0/n515 ), .C0(\U1/aes_core/SB0/n435 ), .C1(
        \U1/aes_core/SB0/n418 ), .Y(\U1/aes_core/SB0/n795 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U471  ( .A(\U1/aes_core/SB0/n400 ), .B(
        \U1/aes_core/SB0/n397 ), .Y(\U1/aes_core/SB0/n635 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U470  ( .A(\U1/aes_core/SB0/n412 ), .B(
        \U1/aes_core/SB0/n491 ), .Y(\U1/aes_core/SB0/n502 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U469  ( .A(\U1/aes_core/SB0/n530 ), .B(
        \U1/aes_core/SB0/n412 ), .Y(\U1/aes_core/SB0/n568 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U468  ( .A(\U1/aes_core/SB0/n546 ), .B(
        \U1/aes_core/SB0/n445 ), .Y(\U1/aes_core/SB0/n696 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U467  ( .AN(\U1/aes_core/SB0/n635 ), .B(
        \U1/aes_core/SB0/n502 ), .C(\U1/aes_core/SB0/n568 ), .D(
        \U1/aes_core/SB0/n696 ), .Y(\U1/aes_core/SB0/n796 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U466  ( .A(\U1/aes_core/SB0/n402 ), .B(
        \U1/aes_core/SB0/n417 ), .Y(\U1/aes_core/SB0/n623 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U465  ( .A(\U1/aes_core/SB0/n546 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n556 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U464  ( .A(\U1/aes_core/SB0/n694 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n655 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U463  ( .A(\U1/aes_core/SB0/n487 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n610 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U462  ( .A(\U1/aes_core/SB0/n623 ), .B(
        \U1/aes_core/SB0/n556 ), .C(\U1/aes_core/SB0/n655 ), .D(
        \U1/aes_core/SB0/n610 ), .Y(\U1/aes_core/SB0/n797 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U461  ( .A(\U1/aes_core/SB0/n794 ), .B(
        \U1/aes_core/SB0/n795 ), .C(\U1/aes_core/SB0/n796 ), .D(
        \U1/aes_core/SB0/n797 ), .Y(\U1/aes_core/SB0/n793 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U460  ( .A(\U1/aes_core/SB0/n793 ), .Y(
        \U1/aes_core/SB0/n420 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U459  ( .A(\U1/aes_core/SB0/n404 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n792 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U458  ( .AN(\U1/aes_core/SB0/n713 ), .B(
        \U1/aes_core/SB0/n791 ), .C(\U1/aes_core/SB0/n420 ), .D(
        \U1/aes_core/SB0/n792 ), .Y(\U1/aes_core/SB0/n790 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U457  ( .A(\U1/aes_core/SB0/n662 ), .B(
        \U1/aes_core/SB0/n565 ), .C(\U1/aes_core/SB0/n787 ), .D(
        \U1/aes_core/SB0/n788 ), .E(\U1/aes_core/SB0/n789 ), .F(
        \U1/aes_core/SB0/n790 ), .Y(\U1/aes_core/SB0/n734 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U456  ( .A(\U1/aes_core/SB0/n419 ), .B(
        \U1/aes_core/SB0/n754 ), .Y(\U1/aes_core/SB0/n617 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U455  ( .A(\U1/aes_core/SB0/n490 ), .B(
        \U1/aes_core/SB0/n402 ), .Y(\U1/aes_core/SB0/n566 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U454  ( .A(\U1/aes_core/SB0/n413 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n664 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U453  ( .A(\U1/aes_core/SB0/n693 ), .Y(
        \U1/aes_core/SB0/n424 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U452  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n641 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U451  ( .AN(\U1/aes_core/SB0/n617 ), .B(
        \U1/aes_core/SB0/n566 ), .C(\U1/aes_core/SB0/n664 ), .D(
        \U1/aes_core/SB0/n641 ), .Y(\U1/aes_core/SB0/n780 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U450  ( .A(\U1/aes_core/SB0/n432 ), .B(
        \U1/aes_core/SB0/n582 ), .Y(\U1/aes_core/SB0/n540 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U449  ( .A(\U1/aes_core/SB0/n530 ), .B(
        \U1/aes_core/SB0/n443 ), .Y(\U1/aes_core/SB0/n684 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U448  ( .A0(\U1/aes_core/SB0/n423 ), .A1(
        \U1/aes_core/SB0/n524 ), .B0(\U1/aes_core/SB0/n694 ), .Y(
        \U1/aes_core/SB0/n786 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U447  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n592 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U446  ( .AN(\U1/aes_core/SB0/n540 ), .B(
        \U1/aes_core/SB0/n684 ), .C(\U1/aes_core/SB0/n786 ), .D(
        \U1/aes_core/SB0/n592 ), .Y(\U1/aes_core/SB0/n785 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U445  ( .A(\U1/aes_core/SB0/n785 ), .Y(
        \U1/aes_core/SB0/n781 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U444  ( .A(\U1/aes_core/SB0/n563 ), .Y(
        \U1/aes_core/SB0/n422 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U443  ( .A(\U1/aes_core/SB0/n397 ), .Y(
        \U1/aes_core/SB0/n523 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U442  ( .A0(\U1/aes_core/SB0/n402 ), 
        .A1(\U1/aes_core/SB0/n489 ), .B0(\U1/aes_core/SB0/n422 ), .B1(
        \U1/aes_core/SB0/n608 ), .C0(\U1/aes_core/SB0/n523 ), .C1(
        \U1/aes_core/SB0/n424 ), .Y(\U1/aes_core/SB0/n782 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U441  ( .A0(\U1/aes_core/SB0/n597 ), .A1(
        \U1/aes_core/SB0/n419 ), .B0(\U1/aes_core/SB0/n399 ), .B1(
        \U1/aes_core/SB0/n398 ), .Y(\U1/aes_core/SB0/n784 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U440  ( .A0(\U1/aes_core/SB0/n546 ), 
        .A1(\U1/aes_core/SB0/n709 ), .B0(\U1/aes_core/SB0/n490 ), .B1(
        \U1/aes_core/SB0/n446 ), .C0(\U1/aes_core/SB0/n784 ), .Y(
        \U1/aes_core/SB0/n783 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U439  ( .AN(\U1/aes_core/SB0/n780 ), .B(
        \U1/aes_core/SB0/n781 ), .C(\U1/aes_core/SB0/n782 ), .D(
        \U1/aes_core/SB0/n783 ), .Y(\U1/aes_core/SB0/n715 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U438  ( .A(\U1/aes_core/SB0/n398 ), .B(
        \U1/aes_core/SB0/n582 ), .Y(\U1/aes_core/SB0/n699 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U437  ( .A0(\U1/aes_core/SB0/n512 ), .A1(
        \U1/aes_core/SB0/n398 ), .B0(\U1/aes_core/SB0/n480 ), .Y(
        \U1/aes_core/SB0/n775 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U436  ( .A(\U1/aes_core/SB0/n480 ), .B(
        \U1/aes_core/SB0/n492 ), .Y(\U1/aes_core/SB0/n615 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB0/U435  ( .A0(\U1/aes_core/SB0/n491 ), .A1(
        \U1/aes_core/SB0/n709 ), .B0(\U1/aes_core/SB0/n615 ), .B1(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n776 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U434  ( .A0(\U1/aes_core/SB0/n437 ), 
        .A1(\U1/aes_core/SB0/n397 ), .B0(\U1/aes_core/SB0/n693 ), .B1(
        \U1/aes_core/SB0/n600 ), .C0(\U1/aes_core/SB0/n435 ), .C1(
        \U1/aes_core/SB0/n406 ), .Y(\U1/aes_core/SB0/n777 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U433  ( .A(\U1/aes_core/SB0/n597 ), .Y(
        \U1/aes_core/SB0/n529 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U432  ( .A(\U1/aes_core/SB0/n404 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n503 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U431  ( .A(\U1/aes_core/SB0/n530 ), .B(
        \U1/aes_core/SB0/n709 ), .Y(\U1/aes_core/SB0/n676 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U430  ( .A(\U1/aes_core/SB0/n694 ), .B(
        \U1/aes_core/SB0/n487 ), .Y(\U1/aes_core/SB0/n656 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U429  ( .A(\U1/aes_core/SB0/n530 ), .B(
        \U1/aes_core/SB0/n489 ), .Y(\U1/aes_core/SB0/n557 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U428  ( .A(\U1/aes_core/SB0/n503 ), .B(
        \U1/aes_core/SB0/n676 ), .C(\U1/aes_core/SB0/n656 ), .D(
        \U1/aes_core/SB0/n557 ), .Y(\U1/aes_core/SB0/n778 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U427  ( .A(\U1/aes_core/SB0/n510 ), .B(
        \U1/aes_core/SB0/n597 ), .Y(\U1/aes_core/SB0/n634 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U426  ( .A(\U1/aes_core/SB0/n524 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n624 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U425  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n608 ), .Y(\U1/aes_core/SB0/n593 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB0/U424  ( .AN(\U1/aes_core/SB0/n634 ), .B(
        \U1/aes_core/SB0/n624 ), .C(\U1/aes_core/SB0/n593 ), .Y(
        \U1/aes_core/SB0/n779 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U423  ( .A(\U1/aes_core/SB0/n699 ), .B(
        \U1/aes_core/SB0/n775 ), .C(\U1/aes_core/SB0/n776 ), .D(
        \U1/aes_core/SB0/n777 ), .E(\U1/aes_core/SB0/n778 ), .F(
        \U1/aes_core/SB0/n779 ), .Y(\U1/aes_core/SB0/n391 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U422  ( .A0(\U1/aes_core/SB0/n694 ), .A1(
        \U1/aes_core/SB0/n445 ), .B0(\U1/aes_core/SB0/n414 ), .Y(
        \U1/aes_core/SB0/n774 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U421  ( .A(\U1/aes_core/SB0/n709 ), .B(
        \U1/aes_core/SB0/n608 ), .Y(\U1/aes_core/SB0/n571 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U420  ( .A(\U1/aes_core/SB0/n491 ), .B(
        \U1/aes_core/SB0/n422 ), .Y(\U1/aes_core/SB0/n679 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U419  ( .A(\U1/aes_core/SB0/n422 ), .B(
        \U1/aes_core/SB0/n487 ), .Y(\U1/aes_core/SB0/n628 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U418  ( .A(\U1/aes_core/SB0/n774 ), .B(
        \U1/aes_core/SB0/n571 ), .C(\U1/aes_core/SB0/n679 ), .D(
        \U1/aes_core/SB0/n628 ), .Y(\U1/aes_core/SB0/n770 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U417  ( .A0(\U1/aes_core/SB0/n419 ), 
        .A1(\U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n693 ), .B1(
        \U1/aes_core/SB0/n447 ), .C0(\U1/aes_core/SB0/n418 ), .C1(
        \U1/aes_core/SB0/n582 ), .Y(\U1/aes_core/SB0/n771 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U416  ( .A(\U1/aes_core/SB0/n488 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n647 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U415  ( .A(\U1/aes_core/SB0/n489 ), .B(
        \U1/aes_core/SB0/n416 ), .Y(\U1/aes_core/SB0/n507 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U414  ( .A(\U1/aes_core/SB0/n489 ), .B(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n660 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U413  ( .A(\U1/aes_core/SB0/n413 ), .B(
        \U1/aes_core/SB0/n423 ), .Y(\U1/aes_core/SB0/n698 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U412  ( .A(\U1/aes_core/SB0/n647 ), .B(
        \U1/aes_core/SB0/n507 ), .C(\U1/aes_core/SB0/n660 ), .D(
        \U1/aes_core/SB0/n698 ), .Y(\U1/aes_core/SB0/n772 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U411  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n585 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U410  ( .A(\U1/aes_core/SB0/n404 ), .B(
        \U1/aes_core/SB0/n443 ), .Y(\U1/aes_core/SB0/n612 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U409  ( .A(\U1/aes_core/SB0/n414 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n561 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U408  ( .A(\U1/aes_core/SB0/n682 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n712 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U407  ( .A(\U1/aes_core/SB0/n585 ), .B(
        \U1/aes_core/SB0/n612 ), .C(\U1/aes_core/SB0/n561 ), .D(
        \U1/aes_core/SB0/n712 ), .Y(\U1/aes_core/SB0/n773 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U406  ( .A(\U1/aes_core/SB0/n770 ), .B(
        \U1/aes_core/SB0/n771 ), .C(\U1/aes_core/SB0/n772 ), .D(
        \U1/aes_core/SB0/n773 ), .Y(\U1/aes_core/SB0/n726 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U405  ( .A(\U1/aes_core/SB0/n734 ), .B(
        \U1/aes_core/SB0/n715 ), .C(\U1/aes_core/SB0/n391 ), .D(
        \U1/aes_core/SB0/n726 ), .Y(\U1/aes_core/SB0/n760 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U404  ( .A(\U1/aes_core/SB0/n437 ), .Y(
        \U1/aes_core/SB0/n534 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U403  ( .A0(\U1/aes_core/SB0/n582 ), .A1(
        \U1/aes_core/SB0/n753 ), .B0(\U1/aes_core/SB0/n613 ), .B1(
        \U1/aes_core/SB0/n406 ), .Y(\U1/aes_core/SB0/n769 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U402  ( .A0(\U1/aes_core/SB0/n534 ), 
        .A1(\U1/aes_core/SB0/n482 ), .B0(\U1/aes_core/SB0/n412 ), .B1(
        \U1/aes_core/SB0/n404 ), .C0(\U1/aes_core/SB0/n769 ), .Y(
        \U1/aes_core/SB0/n761 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U401  ( .A(\U1/aes_core/SB0/n513 ), .B(
        \U1/aes_core/SB0/n510 ), .Y(\U1/aes_core/SB0/n514 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U400  ( .A0(\U1/aes_core/SB0/n579 ), .A1(
        \U1/aes_core/SB0/n510 ), .B0(\U1/aes_core/SB0/n597 ), .B1(
        \U1/aes_core/SB0/n448 ), .Y(\U1/aes_core/SB0/n768 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U399  ( .A0(\U1/aes_core/SB0/n682 ), 
        .A1(\U1/aes_core/SB0/n514 ), .B0(\U1/aes_core/SB0/n442 ), .B1(
        \U1/aes_core/SB0/n423 ), .C0(\U1/aes_core/SB0/n768 ), .Y(
        \U1/aes_core/SB0/n762 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U398  ( .A(\U1/aes_core/SB0/n418 ), .B(
        \U1/aes_core/SB0/n580 ), .Y(\U1/aes_core/SB0/n764 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U397  ( .A(\U1/aes_core/SB0/n489 ), .B(
        \U1/aes_core/SB0/n443 ), .Y(\U1/aes_core/SB0/n522 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U396  ( .A(\U1/aes_core/SB0/n522 ), .Y(
        \U1/aes_core/SB0/n765 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U395  ( .A(\U1/aes_core/SB0/n531 ), .B(
        \U1/aes_core/SB0/n437 ), .Y(\U1/aes_core/SB0/n650 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U394  ( .A(\U1/aes_core/SB0/n432 ), .B(
        \U1/aes_core/SB0/n434 ), .Y(\U1/aes_core/SB0/n497 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U392  ( .A(\U1/aes_core/SB0/n482 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n640 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U390  ( .A0(\U1/aes_core/SB0/n523 ), 
        .A1(\U1/aes_core/SB0/n764 ), .B0(\U1/aes_core/SB0/n546 ), .B1(
        \U1/aes_core/SB0/n765 ), .C0(\U1/aes_core/SB0/n766 ), .Y(
        \U1/aes_core/SB0/n763 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U389  ( .AN(\U1/aes_core/SB0/n760 ), .B(
        \U1/aes_core/SB0/n761 ), .C(\U1/aes_core/SB0/n762 ), .D(
        \U1/aes_core/SB0/n763 ), .Y(\U1/aes_core/sb0 [24]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U388  ( .A(\U1/aes_core/SB0/n510 ), .B(
        \U1/aes_core/SB0/n693 ), .Y(\U1/aes_core/SB0/n633 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U387  ( .A(\U1/aes_core/SB0/n563 ), .B(
        \U1/aes_core/SB0/n513 ), .Y(\U1/aes_core/SB0/n673 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U386  ( .A(\U1/aes_core/SB0/n546 ), .B(
        \U1/aes_core/SB0/n414 ), .Y(\U1/aes_core/SB0/n564 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U385  ( .A0(\U1/aes_core/SB0/n564 ), .A1(
        \U1/aes_core/SB0/n510 ), .B0(\U1/aes_core/SB0/n400 ), .Y(
        \U1/aes_core/SB0/n755 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U384  ( .A(\U1/aes_core/SB0/n482 ), .B(
        \U1/aes_core/SB0/n413 ), .Y(\U1/aes_core/SB0/n657 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U383  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n482 ), .Y(\U1/aes_core/SB0/n558 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U382  ( .A(\U1/aes_core/SB0/n416 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n625 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U381  ( .A(\U1/aes_core/SB0/n657 ), .B(
        \U1/aes_core/SB0/n558 ), .C(\U1/aes_core/SB0/n625 ), .Y(
        \U1/aes_core/SB0/n756 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U380  ( .A(\U1/aes_core/SB0/n482 ), .B(
        \U1/aes_core/SB0/n402 ), .Y(\U1/aes_core/SB0/n598 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U379  ( .A(\U1/aes_core/SB0/n416 ), .B(
        \U1/aes_core/SB0/n425 ), .C(\U1/aes_core/SB0/n404 ), .Y(
        \U1/aes_core/SB0/n759 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U378  ( .A0(\U1/aes_core/SB0/n598 ), 
        .A1(\U1/aes_core/SB0/n436 ), .B0(\U1/aes_core/SB0/n759 ), .B1(
        \U1/aes_core/SB0/n406 ), .C0(\U1/aes_core/SB0/n563 ), .C1(
        \U1/aes_core/SB0/n531 ), .Y(\U1/aes_core/SB0/n757 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U377  ( .A0(\U1/aes_core/SB0/n435 ), .A1(
        \U1/aes_core/SB0/n407 ), .B0(\U1/aes_core/SB0/n434 ), .B1(
        \U1/aes_core/SB0/n437 ), .Y(\U1/aes_core/SB0/n758 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U376  ( .A(\U1/aes_core/SB0/n633 ), .B(
        \U1/aes_core/SB0/n673 ), .C(\U1/aes_core/SB0/n755 ), .D(
        \U1/aes_core/SB0/n756 ), .E(\U1/aes_core/SB0/n757 ), .F(
        \U1/aes_core/SB0/n758 ), .Y(\U1/aes_core/SB0/n392 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U375  ( .A(\U1/aes_core/SB0/n582 ), .B(
        \U1/aes_core/SB0/n597 ), .Y(\U1/aes_core/SB0/n708 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U374  ( .A0(\U1/aes_core/SB0/n582 ), .A1(
        \U1/aes_core/SB0/n492 ), .B0(\U1/aes_core/SB0/n693 ), .Y(
        \U1/aes_core/SB0/n747 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U373  ( .A(\U1/aes_core/SB0/n488 ), .B(
        \U1/aes_core/SB0/n482 ), .Y(\U1/aes_core/SB0/n705 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U372  ( .A0(\U1/aes_core/SB0/n600 ), .A1(
        \U1/aes_core/SB0/n432 ), .B0(\U1/aes_core/SB0/n705 ), .B1(
        \U1/aes_core/SB0/n418 ), .Y(\U1/aes_core/SB0/n748 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U371  ( .A0(\U1/aes_core/SB0/n613 ), 
        .A1(\U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n448 ), .B1(
        \U1/aes_core/SB0/n563 ), .C0(\U1/aes_core/SB0/n434 ), .C1(
        \U1/aes_core/SB0/n512 ), .Y(\U1/aes_core/SB0/n749 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U370  ( .A(\U1/aes_core/SB0/n399 ), .B(
        \U1/aes_core/SB0/n754 ), .Y(\U1/aes_core/SB0/n649 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U369  ( .A(\U1/aes_core/SB0/n412 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n642 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U368  ( .A(\U1/aes_core/SB0/n491 ), .B(
        \U1/aes_core/SB0/n417 ), .Y(\U1/aes_core/SB0/n632 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U367  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n402 ), .Y(\U1/aes_core/SB0/n528 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U366  ( .AN(\U1/aes_core/SB0/n649 ), .B(
        \U1/aes_core/SB0/n642 ), .C(\U1/aes_core/SB0/n632 ), .D(
        \U1/aes_core/SB0/n528 ), .Y(\U1/aes_core/SB0/n750 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U365  ( .A(\U1/aes_core/SB0/n531 ), .B(
        \U1/aes_core/SB0/n753 ), .Y(\U1/aes_core/SB0/n549 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U364  ( .A(\U1/aes_core/SB0/n432 ), .B(
        \U1/aes_core/SB0/n448 ), .Y(\U1/aes_core/SB0/n496 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U362  ( .A(\U1/aes_core/SB0/n709 ), .B(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n683 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U360  ( .A(\U1/aes_core/SB0/n708 ), .B(
        \U1/aes_core/SB0/n747 ), .C(\U1/aes_core/SB0/n748 ), .D(
        \U1/aes_core/SB0/n749 ), .E(\U1/aes_core/SB0/n750 ), .F(
        \U1/aes_core/SB0/n751 ), .Y(\U1/aes_core/SB0/n714 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U359  ( .A(\U1/aes_core/SB0/n515 ), .B(
        \U1/aes_core/SB0/n693 ), .Y(\U1/aes_core/SB0/n695 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U358  ( .A(\U1/aes_core/SB0/n563 ), .B(
        \U1/aes_core/SB0/n613 ), .Y(\U1/aes_core/SB0/n483 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U357  ( .A(\U1/aes_core/SB0/n582 ), .B(
        \U1/aes_core/SB0/n512 ), .Y(\U1/aes_core/SB0/n645 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U356  ( .A(\U1/aes_core/SB0/n397 ), .B(
        \U1/aes_core/SB0/n512 ), .Y(\U1/aes_core/SB0/n630 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U355  ( .A(\U1/aes_core/SB0/n487 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n570 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U354  ( .A(\U1/aes_core/SB0/n416 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n678 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U353  ( .A(\U1/aes_core/SB0/n412 ), .B(
        \U1/aes_core/SB0/n416 ), .Y(\U1/aes_core/SB0/n584 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U352  ( .A(\U1/aes_core/SB0/n523 ), .B(
        \U1/aes_core/SB0/n445 ), .Y(\U1/aes_core/SB0/n659 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U351  ( .A(\U1/aes_core/SB0/n570 ), .B(
        \U1/aes_core/SB0/n678 ), .C(\U1/aes_core/SB0/n584 ), .D(
        \U1/aes_core/SB0/n659 ), .Y(\U1/aes_core/SB0/n743 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U350  ( .A(\U1/aes_core/SB0/n397 ), .B(
        \U1/aes_core/SB0/n597 ), .Y(\U1/aes_core/SB0/n609 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U349  ( .A(\U1/aes_core/SB0/n398 ), .B(
        \U1/aes_core/SB0/n613 ), .Y(\U1/aes_core/SB0/n509 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U348  ( .A(\U1/aes_core/SB0/n492 ), .B(
        \U1/aes_core/SB0/n432 ), .Y(\U1/aes_core/SB0/n559 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U347  ( .A(\U1/aes_core/SB0/n531 ), .B(
        \U1/aes_core/SB0/n432 ), .Y(\U1/aes_core/SB0/n710 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U346  ( .A0(\U1/aes_core/SB0/n432 ), .A1(
        \U1/aes_core/SB0/n397 ), .B0(\U1/aes_core/SB0/n597 ), .B1(
        \U1/aes_core/SB0/n492 ), .Y(\U1/aes_core/SB0/n745 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U345  ( .A0(\U1/aes_core/SB0/n613 ), .A1(
        \U1/aes_core/SB0/n400 ), .B0(\U1/aes_core/SB0/n600 ), .B1(
        \U1/aes_core/SB0/n563 ), .Y(\U1/aes_core/SB0/n746 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U344  ( .A(\U1/aes_core/SB0/n609 ), .B(
        \U1/aes_core/SB0/n509 ), .C(\U1/aes_core/SB0/n559 ), .D(
        \U1/aes_core/SB0/n710 ), .E(\U1/aes_core/SB0/n745 ), .F(
        \U1/aes_core/SB0/n746 ), .Y(\U1/aes_core/SB0/n744 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U343  ( .A(\U1/aes_core/SB0/n695 ), .B(
        \U1/aes_core/SB0/n483 ), .C(\U1/aes_core/SB0/n645 ), .D(
        \U1/aes_core/SB0/n630 ), .E(\U1/aes_core/SB0/n743 ), .F(
        \U1/aes_core/SB0/n744 ), .Y(\U1/aes_core/SB0/n725 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U342  ( .A0(\U1/aes_core/SB0/n487 ), 
        .A1(\U1/aes_core/SB0/n490 ), .B0(\U1/aes_core/SB0/n413 ), .B1(
        \U1/aes_core/SB0/n546 ), .C0(\U1/aes_core/SB0/n725 ), .Y(
        \U1/aes_core/SB0/n742 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U341  ( .A(\U1/aes_core/SB0/n742 ), .Y(
        \U1/aes_core/SB0/n735 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U340  ( .A(\U1/aes_core/SB0/n434 ), .B(
        \U1/aes_core/SB0/n492 ), .Y(\U1/aes_core/SB0/n444 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U339  ( .A0(\U1/aes_core/SB0/n488 ), .A1(
        \U1/aes_core/SB0/n444 ), .B0(\U1/aes_core/SB0/n412 ), .Y(
        \U1/aes_core/SB0/n739 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U338  ( .A0(\U1/aes_core/SB0/n523 ), .A1(
        \U1/aes_core/SB0/n423 ), .B0(\U1/aes_core/SB0/n481 ), .Y(
        \U1/aes_core/SB0/n740 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U337  ( .A0(\U1/aes_core/SB0/n524 ), .A1(
        \U1/aes_core/SB0/n482 ), .B0(\U1/aes_core/SB0/n417 ), .Y(
        \U1/aes_core/SB0/n741 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U336  ( .A(\U1/aes_core/SB0/n491 ), .B(
        \U1/aes_core/SB0/n424 ), .Y(\U1/aes_core/SB0/n666 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U335  ( .A(\U1/aes_core/SB0/n739 ), .B(
        \U1/aes_core/SB0/n740 ), .C(\U1/aes_core/SB0/n741 ), .D(
        \U1/aes_core/SB0/n666 ), .Y(\U1/aes_core/SB0/n736 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U334  ( .A(\U1/aes_core/SB0/n425 ), .B(
        \U1/aes_core/SB0/n530 ), .Y(\U1/aes_core/SB0/n476 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB0/U333  ( .A(\U1/aes_core/SB0/n476 ), .B(
        \U1/aes_core/SB0/n435 ), .C(\U1/aes_core/SB0/n448 ), .Y(
        \U1/aes_core/SB0/n738 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U332  ( .A0(\U1/aes_core/SB0/n492 ), 
        .A1(\U1/aes_core/SB0/n398 ), .B0(\U1/aes_core/SB0/n738 ), .B1(
        \U1/aes_core/SB0/n437 ), .C0(\U1/aes_core/SB0/n399 ), .C1(
        \U1/aes_core/SB0/n407 ), .Y(\U1/aes_core/SB0/n737 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U331  ( .A(\U1/aes_core/SB0/n392 ), .B(
        \U1/aes_core/SB0/n714 ), .C(\U1/aes_core/SB0/n734 ), .D(
        \U1/aes_core/SB0/n735 ), .E(\U1/aes_core/SB0/n736 ), .F(
        \U1/aes_core/SB0/n737 ), .Y(\U1/aes_core/sb0 [25]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U330  ( .A0(\U1/aes_core/SB0/n443 ), .A1(
        \U1/aes_core/SB0/n423 ), .B0(\U1/aes_core/SB0/n402 ), .B1(
        \U1/aes_core/SB0/n412 ), .Y(\U1/aes_core/SB0/n733 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U329  ( .A0(\U1/aes_core/SB0/n513 ), 
        .A1(\U1/aes_core/SB0/n398 ), .B0(\U1/aes_core/SB0/n563 ), .B1(
        \U1/aes_core/SB0/n492 ), .C0(\U1/aes_core/SB0/n733 ), .Y(
        \U1/aes_core/SB0/n727 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U328  ( .A(\U1/aes_core/SB0/n417 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n629 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U327  ( .A(\U1/aes_core/SB0/n443 ), .B(
        \U1/aes_core/SB0/n488 ), .Y(\U1/aes_core/SB0/n648 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U326  ( .A(\U1/aes_core/SB0/n423 ), .B(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n680 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U325  ( .A(\U1/aes_core/SB0/n524 ), .B(
        \U1/aes_core/SB0/n481 ), .Y(\U1/aes_core/SB0/n661 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U324  ( .A(\U1/aes_core/SB0/n629 ), .B(
        \U1/aes_core/SB0/n648 ), .C(\U1/aes_core/SB0/n680 ), .D(
        \U1/aes_core/SB0/n661 ), .Y(\U1/aes_core/SB0/n728 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U323  ( .A(\U1/aes_core/SB0/n397 ), .B(
        \U1/aes_core/SB0/n419 ), .Y(\U1/aes_core/SB0/n535 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U322  ( .A0(\U1/aes_core/SB0/n487 ), .A1(
        \U1/aes_core/SB0/n535 ), .B0(\U1/aes_core/SB0/n413 ), .Y(
        \U1/aes_core/SB0/n730 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U321  ( .A0(\U1/aes_core/SB0/n416 ), .A1(
        \U1/aes_core/SB0/n546 ), .B0(\U1/aes_core/SB0/n534 ), .Y(
        \U1/aes_core/SB0/n731 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U320  ( .A0(\U1/aes_core/SB0/n529 ), .A1(
        \U1/aes_core/SB0/n489 ), .B0(\U1/aes_core/SB0/n414 ), .Y(
        \U1/aes_core/SB0/n732 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U319  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n416 ), .Y(\U1/aes_core/SB0/n562 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U318  ( .A(\U1/aes_core/SB0/n730 ), .B(
        \U1/aes_core/SB0/n731 ), .C(\U1/aes_core/SB0/n732 ), .D(
        \U1/aes_core/SB0/n562 ), .Y(\U1/aes_core/SB0/n729 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U317  ( .A(\U1/aes_core/SB0/n724 ), .B(
        \U1/aes_core/SB0/n725 ), .C(\U1/aes_core/SB0/n726 ), .D(
        \U1/aes_core/SB0/n727 ), .E(\U1/aes_core/SB0/n728 ), .F(
        \U1/aes_core/SB0/n729 ), .Y(\U1/aes_core/SB0/n393 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U316  ( .A0(\U1/aes_core/SB0/n608 ), 
        .A1(\U1/aes_core/SB0/n412 ), .B0(\U1/aes_core/SB0/n404 ), .B1(
        \U1/aes_core/SB0/n490 ), .C0(\U1/aes_core/SB0/n393 ), .Y(
        \U1/aes_core/SB0/n723 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U315  ( .A(\U1/aes_core/SB0/n723 ), .Y(
        \U1/aes_core/SB0/n716 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U314  ( .A(\U1/aes_core/SB0/n481 ), .B(
        \U1/aes_core/SB0/n694 ), .Y(\U1/aes_core/SB0/n572 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U313  ( .A1N(\U1/aes_core/SB0/n572 ), 
        .A0(\U1/aes_core/SB0/n442 ), .B0(\U1/aes_core/SB0/n491 ), .Y(
        \U1/aes_core/SB0/n720 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U312  ( .A0(\U1/aes_core/SB0/n523 ), .A1(
        \U1/aes_core/SB0/n615 ), .B0(\U1/aes_core/SB0/n443 ), .Y(
        \U1/aes_core/SB0/n721 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U311  ( .A0(\U1/aes_core/SB0/n416 ), .A1(
        \U1/aes_core/SB0/n482 ), .B0(\U1/aes_core/SB0/n422 ), .Y(
        \U1/aes_core/SB0/n722 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U310  ( .A(\U1/aes_core/SB0/n445 ), .B(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n665 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U309  ( .A(\U1/aes_core/SB0/n720 ), .B(
        \U1/aes_core/SB0/n721 ), .C(\U1/aes_core/SB0/n722 ), .D(
        \U1/aes_core/SB0/n665 ), .Y(\U1/aes_core/SB0/n717 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U308  ( .A(\U1/aes_core/SB0/n446 ), .B(
        \U1/aes_core/SB0/n414 ), .Y(\U1/aes_core/SB0/n415 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U307  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n489 ), .Y(\U1/aes_core/SB0/n719 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U306  ( .A0(\U1/aes_core/SB0/n415 ), 
        .A1(\U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n719 ), .B1(
        \U1/aes_core/SB0/n434 ), .C0(\U1/aes_core/SB0/n512 ), .C1(
        \U1/aes_core/SB0/n510 ), .Y(\U1/aes_core/SB0/n718 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U305  ( .A(\U1/aes_core/SB0/n713 ), .B(
        \U1/aes_core/SB0/n714 ), .C(\U1/aes_core/SB0/n715 ), .D(
        \U1/aes_core/SB0/n716 ), .E(\U1/aes_core/SB0/n717 ), .F(
        \U1/aes_core/SB0/n718 ), .Y(\U1/aes_core/sb0 [26]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U304  ( .A(\U1/aes_core/SB0/n608 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n410 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U303  ( .AN(\U1/aes_core/SB0/n710 ), .B(
        \U1/aes_core/SB0/n711 ), .C(\U1/aes_core/SB0/n712 ), .D(
        \U1/aes_core/SB0/n410 ), .Y(\U1/aes_core/SB0/n702 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U302  ( .A0(\U1/aes_core/SB0/n709 ), .A1(
        \U1/aes_core/SB0/n443 ), .B0(\U1/aes_core/SB0/n546 ), .Y(
        \U1/aes_core/SB0/n706 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U299  ( .A(\U1/aes_core/SB0/n490 ), .B(
        \U1/aes_core/SB0/n422 ), .Y(\U1/aes_core/SB0/n479 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U298  ( .A0(\U1/aes_core/SB0/n600 ), 
        .A1(\U1/aes_core/SB0/n400 ), .B0(\U1/aes_core/SB0/n479 ), .B1(
        \U1/aes_core/SB0/n447 ), .C0(\U1/aes_core/SB0/n406 ), .C1(
        \U1/aes_core/SB0/n397 ), .Y(\U1/aes_core/SB0/n704 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U297  ( .A(\U1/aes_core/SB0/n699 ), .B(
        \U1/aes_core/SB0/n700 ), .C(\U1/aes_core/SB0/n701 ), .D(
        \U1/aes_core/SB0/n702 ), .E(\U1/aes_core/SB0/n703 ), .F(
        \U1/aes_core/SB0/n704 ), .Y(\U1/aes_core/SB0/n516 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U296  ( .AN(\U1/aes_core/SB0/n695 ), .B(
        \U1/aes_core/SB0/n696 ), .C(\U1/aes_core/SB0/n697 ), .D(
        \U1/aes_core/SB0/n698 ), .Y(\U1/aes_core/SB0/n685 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U295  ( .A0(\U1/aes_core/SB0/n412 ), 
        .A1(\U1/aes_core/SB0/n523 ), .B0(\U1/aes_core/SB0/n417 ), .B1(
        \U1/aes_core/SB0/n524 ), .C0(\U1/aes_core/SB0/n694 ), .C1(
        \U1/aes_core/SB0/n402 ), .Y(\U1/aes_core/SB0/n686 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U294  ( .A0(\U1/aes_core/SB0/n448 ), .A1(
        \U1/aes_core/SB0/n563 ), .B0(\U1/aes_core/SB0/n693 ), .B1(
        \U1/aes_core/SB0/n600 ), .Y(\U1/aes_core/SB0/n692 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U293  ( .A0(\U1/aes_core/SB0/n546 ), 
        .A1(\U1/aes_core/SB0/n529 ), .B0(\U1/aes_core/SB0/n530 ), .B1(
        \U1/aes_core/SB0/n445 ), .C0(\U1/aes_core/SB0/n692 ), .Y(
        \U1/aes_core/SB0/n687 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U292  ( .A(\U1/aes_core/SB0/n437 ), .B(
        \U1/aes_core/SB0/n398 ), .Y(\U1/aes_core/SB0/n690 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U291  ( .A0(\U1/aes_core/SB0/n608 ), 
        .A1(\U1/aes_core/SB0/n689 ), .B0(\U1/aes_core/SB0/n416 ), .B1(
        \U1/aes_core/SB0/n690 ), .C0(\U1/aes_core/SB0/n691 ), .Y(
        \U1/aes_core/SB0/n688 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U290  ( .AN(\U1/aes_core/SB0/n685 ), .B(
        \U1/aes_core/SB0/n686 ), .C(\U1/aes_core/SB0/n687 ), .D(
        \U1/aes_core/SB0/n688 ), .Y(\U1/aes_core/SB0/n471 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U289  ( .A(\U1/aes_core/SB0/n684 ), .Y(
        \U1/aes_core/SB0/n668 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U288  ( .A0(\U1/aes_core/SB0/n579 ), .A1(
        \U1/aes_core/SB0/n510 ), .B0(\U1/aes_core/SB0/n683 ), .Y(
        \U1/aes_core/SB0/n669 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U287  ( .A0(\U1/aes_core/SB0/n416 ), .A1(
        \U1/aes_core/SB0/n417 ), .B0(\U1/aes_core/SB0/n446 ), .B1(
        \U1/aes_core/SB0/n682 ), .Y(\U1/aes_core/SB0/n681 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U286  ( .A0(\U1/aes_core/SB0/n435 ), 
        .A1(\U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n419 ), .B1(
        \U1/aes_core/SB0/n407 ), .C0(\U1/aes_core/SB0/n681 ), .Y(
        \U1/aes_core/SB0/n670 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U285  ( .A(\U1/aes_core/SB0/n677 ), .B(
        \U1/aes_core/SB0/n678 ), .C(\U1/aes_core/SB0/n679 ), .D(
        \U1/aes_core/SB0/n680 ), .Y(\U1/aes_core/SB0/n671 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U284  ( .AN(\U1/aes_core/SB0/n673 ), .B(
        \U1/aes_core/SB0/n674 ), .C(\U1/aes_core/SB0/n675 ), .D(
        \U1/aes_core/SB0/n676 ), .Y(\U1/aes_core/SB0/n672 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U283  ( .A(\U1/aes_core/SB0/n667 ), .B(
        \U1/aes_core/SB0/n668 ), .C(\U1/aes_core/SB0/n669 ), .D(
        \U1/aes_core/SB0/n670 ), .E(\U1/aes_core/SB0/n671 ), .F(
        \U1/aes_core/SB0/n672 ), .Y(\U1/aes_core/SB0/n567 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U282  ( .A0(\U1/aes_core/SB0/n480 ), .A1(
        \U1/aes_core/SB0/n563 ), .B0(\U1/aes_core/SB0/n666 ), .Y(
        \U1/aes_core/SB0/n651 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U281  ( .AN(\U1/aes_core/SB0/n662 ), .B(
        \U1/aes_core/SB0/n663 ), .C(\U1/aes_core/SB0/n664 ), .D(
        \U1/aes_core/SB0/n665 ), .Y(\U1/aes_core/SB0/n652 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U280  ( .A(\U1/aes_core/SB0/n425 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n411 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U279  ( .A(\U1/aes_core/SB0/n659 ), .B(
        \U1/aes_core/SB0/n660 ), .C(\U1/aes_core/SB0/n661 ), .D(
        \U1/aes_core/SB0/n411 ), .Y(\U1/aes_core/SB0/n653 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U278  ( .A(\U1/aes_core/SB0/n655 ), .B(
        \U1/aes_core/SB0/n656 ), .C(\U1/aes_core/SB0/n657 ), .D(
        \U1/aes_core/SB0/n658 ), .Y(\U1/aes_core/SB0/n654 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U277  ( .A(\U1/aes_core/SB0/n649 ), .B(
        \U1/aes_core/SB0/n650 ), .C(\U1/aes_core/SB0/n651 ), .D(
        \U1/aes_core/SB0/n652 ), .E(\U1/aes_core/SB0/n653 ), .F(
        \U1/aes_core/SB0/n654 ), .Y(\U1/aes_core/SB0/n543 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U276  ( .AN(\U1/aes_core/SB0/n645 ), .B(
        \U1/aes_core/SB0/n646 ), .C(\U1/aes_core/SB0/n647 ), .D(
        \U1/aes_core/SB0/n648 ), .Y(\U1/aes_core/SB0/n636 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U275  ( .A(\U1/aes_core/SB0/n641 ), .B(
        \U1/aes_core/SB0/n642 ), .C(\U1/aes_core/SB0/n643 ), .D(
        \U1/aes_core/SB0/n644 ), .Y(\U1/aes_core/SB0/n637 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U274  ( .A(\U1/aes_core/SB0/n481 ), .B(
        \U1/aes_core/SB0/n424 ), .C(\U1/aes_core/SB0/n422 ), .Y(
        \U1/aes_core/SB0/n639 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U273  ( .A0(\U1/aes_core/SB0/n639 ), 
        .A1(\U1/aes_core/SB0/n434 ), .B0(\U1/aes_core/SB0/n600 ), .B1(
        \U1/aes_core/SB0/n398 ), .C0(\U1/aes_core/SB0/n640 ), .Y(
        \U1/aes_core/SB0/n638 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U272  ( .A(\U1/aes_core/SB0/n633 ), .B(
        \U1/aes_core/SB0/n634 ), .C(\U1/aes_core/SB0/n635 ), .D(
        \U1/aes_core/SB0/n636 ), .E(\U1/aes_core/SB0/n637 ), .F(
        \U1/aes_core/SB0/n638 ), .Y(\U1/aes_core/SB0/n495 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U271  ( .A0(\U1/aes_core/SB0/n600 ), .A1(
        \U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n632 ), .Y(
        \U1/aes_core/SB0/n618 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U270  ( .A0(\U1/aes_core/SB0/n491 ), .A1(
        \U1/aes_core/SB0/n489 ), .B0(\U1/aes_core/SB0/n413 ), .B1(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n631 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U269  ( .A0(\U1/aes_core/SB0/n580 ), 
        .A1(\U1/aes_core/SB0/n492 ), .B0(\U1/aes_core/SB0/n579 ), .B1(
        \U1/aes_core/SB0/n515 ), .C0(\U1/aes_core/SB0/n631 ), .Y(
        \U1/aes_core/SB0/n619 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U268  ( .A(\U1/aes_core/SB0/n630 ), .Y(
        \U1/aes_core/SB0/n627 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U267  ( .AN(\U1/aes_core/SB0/n626 ), .B(
        \U1/aes_core/SB0/n627 ), .C(\U1/aes_core/SB0/n628 ), .D(
        \U1/aes_core/SB0/n629 ), .Y(\U1/aes_core/SB0/n620 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U266  ( .A(\U1/aes_core/SB0/n622 ), .B(
        \U1/aes_core/SB0/n623 ), .C(\U1/aes_core/SB0/n624 ), .D(
        \U1/aes_core/SB0/n625 ), .Y(\U1/aes_core/SB0/n621 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U265  ( .A(\U1/aes_core/SB0/n616 ), .B(
        \U1/aes_core/SB0/n617 ), .C(\U1/aes_core/SB0/n618 ), .D(
        \U1/aes_core/SB0/n619 ), .E(\U1/aes_core/SB0/n620 ), .F(
        \U1/aes_core/SB0/n621 ), .Y(\U1/aes_core/SB0/n536 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U264  ( .A0(\U1/aes_core/SB0/n424 ), .A1(
        \U1/aes_core/SB0/n615 ), .B0(\U1/aes_core/SB0/n414 ), .B1(
        \U1/aes_core/SB0/n489 ), .Y(\U1/aes_core/SB0/n614 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U263  ( .A0(\U1/aes_core/SB0/n563 ), 
        .A1(\U1/aes_core/SB0/n397 ), .B0(\U1/aes_core/SB0/n613 ), .B1(
        \U1/aes_core/SB0/n407 ), .C0(\U1/aes_core/SB0/n614 ), .Y(
        \U1/aes_core/SB0/n601 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U262  ( .AN(\U1/aes_core/SB0/n609 ), .B(
        \U1/aes_core/SB0/n610 ), .C(\U1/aes_core/SB0/n611 ), .D(
        \U1/aes_core/SB0/n612 ), .Y(\U1/aes_core/SB0/n602 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U261  ( .A0(\U1/aes_core/SB0/n404 ), .A1(
        \U1/aes_core/SB0/n608 ), .B0(\U1/aes_core/SB0/n413 ), .Y(
        \U1/aes_core/SB0/n604 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U260  ( .A(\U1/aes_core/SB0/n437 ), .B(
        \U1/aes_core/SB0/n432 ), .Y(\U1/aes_core/SB0/n607 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U259  ( .A0(\U1/aes_core/SB0/n482 ), .A1(
        \U1/aes_core/SB0/n607 ), .B0(\U1/aes_core/SB0/n481 ), .B1(
        \U1/aes_core/SB0/n535 ), .Y(\U1/aes_core/SB0/n606 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U258  ( .A(\U1/aes_core/SB0/n604 ), .B(
        \U1/aes_core/SB0/n605 ), .C(\U1/aes_core/SB0/n606 ), .Y(
        \U1/aes_core/SB0/n603 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U257  ( .A(\U1/aes_core/SB0/n543 ), .B(
        \U1/aes_core/SB0/n495 ), .C(\U1/aes_core/SB0/n536 ), .D(
        \U1/aes_core/SB0/n601 ), .E(\U1/aes_core/SB0/n602 ), .F(
        \U1/aes_core/SB0/n603 ), .Y(\U1/aes_core/SB0/n428 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U256  ( .A(\U1/aes_core/SB0/n516 ), .B(
        \U1/aes_core/SB0/n471 ), .C(\U1/aes_core/SB0/n567 ), .D(
        \U1/aes_core/SB0/n428 ), .Y(\U1/aes_core/SB0/n587 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U255  ( .A0(\U1/aes_core/SB0/n448 ), .A1(
        \U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n600 ), .B1(
        \U1/aes_core/SB0/n432 ), .Y(\U1/aes_core/SB0/n599 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U254  ( .A0(\U1/aes_core/SB0/n443 ), 
        .A1(\U1/aes_core/SB0/n425 ), .B0(\U1/aes_core/SB0/n412 ), .B1(
        \U1/aes_core/SB0/n404 ), .C0(\U1/aes_core/SB0/n599 ), .Y(
        \U1/aes_core/SB0/n588 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U253  ( .A(\U1/aes_core/SB0/n598 ), .Y(
        \U1/aes_core/SB0/n595 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U252  ( .A0(\U1/aes_core/SB0/n597 ), .A1(
        \U1/aes_core/SB0/n492 ), .B0(\U1/aes_core/SB0/n564 ), .B1(
        \U1/aes_core/SB0/n512 ), .Y(\U1/aes_core/SB0/n596 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U251  ( .A0(\U1/aes_core/SB0/n424 ), 
        .A1(\U1/aes_core/SB0/n595 ), .B0(\U1/aes_core/SB0/n442 ), .B1(
        \U1/aes_core/SB0/n514 ), .C0(\U1/aes_core/SB0/n596 ), .Y(
        \U1/aes_core/SB0/n589 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U250  ( .A0(\U1/aes_core/SB0/n402 ), .A1(
        \U1/aes_core/SB0/n546 ), .B0(\U1/aes_core/SB0/n422 ), .Y(
        \U1/aes_core/SB0/n591 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB0/U249  ( .A(\U1/aes_core/SB0/n591 ), .B(
        \U1/aes_core/SB0/n592 ), .C(\U1/aes_core/SB0/n593 ), .D(
        \U1/aes_core/SB0/n594 ), .Y(\U1/aes_core/SB0/n590 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U248  ( .AN(\U1/aes_core/SB0/n587 ), .B(
        \U1/aes_core/SB0/n588 ), .C(\U1/aes_core/SB0/n589 ), .D(
        \U1/aes_core/SB0/n590 ), .Y(\U1/aes_core/sb0 [27]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U247  ( .A0(\U1/aes_core/SB0/n572 ), .A1(
        \U1/aes_core/SB0/n436 ), .B0(\U1/aes_core/SB0/n513 ), .Y(
        \U1/aes_core/SB0/n575 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U246  ( .A(\U1/aes_core/SB0/n584 ), .B(
        \U1/aes_core/SB0/n585 ), .C(\U1/aes_core/SB0/n586 ), .Y(
        \U1/aes_core/SB0/n576 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U245  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n413 ), .Y(\U1/aes_core/SB0/n581 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U244  ( .A(\U1/aes_core/SB0/n442 ), .B(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n583 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U243  ( .A0(\U1/aes_core/SB0/n581 ), 
        .A1(\U1/aes_core/SB0/n582 ), .B0(\U1/aes_core/SB0/n583 ), .B1(
        \U1/aes_core/SB0/n419 ), .C0(\U1/aes_core/SB0/n436 ), .C1(
        \U1/aes_core/SB0/n531 ), .Y(\U1/aes_core/SB0/n577 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U242  ( .A0(\U1/aes_core/SB0/n480 ), 
        .A1(\U1/aes_core/SB0/n579 ), .B0(\U1/aes_core/SB0/n397 ), .B1(
        \U1/aes_core/SB0/n407 ), .C0(\U1/aes_core/SB0/n434 ), .C1(
        \U1/aes_core/SB0/n580 ), .Y(\U1/aes_core/SB0/n578 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U241  ( .A(\U1/aes_core/SB0/n573 ), .B(
        \U1/aes_core/SB0/n574 ), .C(\U1/aes_core/SB0/n575 ), .D(
        \U1/aes_core/SB0/n576 ), .E(\U1/aes_core/SB0/n577 ), .F(
        \U1/aes_core/SB0/n578 ), .Y(\U1/aes_core/SB0/n427 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U240  ( .A0(\U1/aes_core/SB0/n572 ), .A1(
        \U1/aes_core/SB0/n563 ), .B0(\U1/aes_core/SB0/n492 ), .Y(
        \U1/aes_core/SB0/n537 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB0/U239  ( .A0(\U1/aes_core/SB0/n447 ), .A1(
        \U1/aes_core/SB0/n434 ), .A2(\U1/aes_core/SB0/n515 ), .B0(
        \U1/aes_core/SB0/n418 ), .Y(\U1/aes_core/SB0/n538 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U238  ( .A(\U1/aes_core/SB0/n568 ), .B(
        \U1/aes_core/SB0/n569 ), .C(\U1/aes_core/SB0/n570 ), .D(
        \U1/aes_core/SB0/n571 ), .Y(\U1/aes_core/SB0/n541 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U237  ( .A(\U1/aes_core/SB0/n567 ), .Y(
        \U1/aes_core/SB0/n544 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U236  ( .A(\U1/aes_core/SB0/n566 ), .Y(
        \U1/aes_core/SB0/n550 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB0/U235  ( .A0(\U1/aes_core/SB0/n564 ), 
        .A1(\U1/aes_core/SB0/n406 ), .B0N(\U1/aes_core/SB0/n565 ), .Y(
        \U1/aes_core/SB0/n551 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U234  ( .A0(\U1/aes_core/SB0/n399 ), 
        .A1(\U1/aes_core/SB0/n563 ), .B0(\U1/aes_core/SB0/n513 ), .B1(
        \U1/aes_core/SB0/n432 ), .C0(\U1/aes_core/SB0/n418 ), .C1(
        \U1/aes_core/SB0/n397 ), .Y(\U1/aes_core/SB0/n552 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U233  ( .AN(\U1/aes_core/SB0/n559 ), .B(
        \U1/aes_core/SB0/n560 ), .C(\U1/aes_core/SB0/n561 ), .D(
        \U1/aes_core/SB0/n562 ), .Y(\U1/aes_core/SB0/n553 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U232  ( .A(\U1/aes_core/SB0/n555 ), .B(
        \U1/aes_core/SB0/n556 ), .C(\U1/aes_core/SB0/n557 ), .D(
        \U1/aes_core/SB0/n558 ), .Y(\U1/aes_core/SB0/n554 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U231  ( .A(\U1/aes_core/SB0/n549 ), .B(
        \U1/aes_core/SB0/n550 ), .C(\U1/aes_core/SB0/n551 ), .D(
        \U1/aes_core/SB0/n552 ), .E(\U1/aes_core/SB0/n553 ), .F(
        \U1/aes_core/SB0/n554 ), .Y(\U1/aes_core/SB0/n548 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U230  ( .A(\U1/aes_core/SB0/n548 ), .Y(
        \U1/aes_core/SB0/n449 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U229  ( .A0(\U1/aes_core/SB0/n480 ), .A1(
        \U1/aes_core/SB0/n437 ), .B0(\U1/aes_core/SB0/n397 ), .B1(
        \U1/aes_core/SB0/n398 ), .Y(\U1/aes_core/SB0/n547 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U228  ( .A0(\U1/aes_core/SB0/n490 ), 
        .A1(\U1/aes_core/SB0/n546 ), .B0(\U1/aes_core/SB0/n445 ), .B1(
        \U1/aes_core/SB0/n423 ), .C0(\U1/aes_core/SB0/n547 ), .Y(
        \U1/aes_core/SB0/n545 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U227  ( .AN(\U1/aes_core/SB0/n543 ), .B(
        \U1/aes_core/SB0/n544 ), .C(\U1/aes_core/SB0/n449 ), .D(
        \U1/aes_core/SB0/n545 ), .Y(\U1/aes_core/SB0/n542 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U226  ( .A(\U1/aes_core/SB0/n537 ), .B(
        \U1/aes_core/SB0/n538 ), .C(\U1/aes_core/SB0/n539 ), .D(
        \U1/aes_core/SB0/n540 ), .E(\U1/aes_core/SB0/n541 ), .F(
        \U1/aes_core/SB0/n542 ), .Y(\U1/aes_core/SB0/n472 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U225  ( .A(\U1/aes_core/SB0/n536 ), .Y(
        \U1/aes_core/SB0/n532 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U224  ( .A0(\U1/aes_core/SB0/n534 ), .A1(
        \U1/aes_core/SB0/n535 ), .B0(\U1/aes_core/SB0/n488 ), .B1(
        \U1/aes_core/SB0/n529 ), .Y(\U1/aes_core/SB0/n533 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U223  ( .A0(\U1/aes_core/SB0/n418 ), 
        .A1(\U1/aes_core/SB0/n531 ), .B0(\U1/aes_core/SB0/n532 ), .C0(
        \U1/aes_core/SB0/n533 ), .Y(\U1/aes_core/SB0/n517 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U222  ( .A0(\U1/aes_core/SB0/n530 ), .A1(
        \U1/aes_core/SB0/n446 ), .B0(\U1/aes_core/SB0/n417 ), .Y(
        \U1/aes_core/SB0/n525 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U221  ( .A0(\U1/aes_core/SB0/n529 ), .A1(
        \U1/aes_core/SB0/n443 ), .B0(\U1/aes_core/SB0/n414 ), .Y(
        \U1/aes_core/SB0/n526 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U220  ( .A(\U1/aes_core/SB0/n525 ), .B(
        \U1/aes_core/SB0/n526 ), .C(\U1/aes_core/SB0/n527 ), .D(
        \U1/aes_core/SB0/n528 ), .Y(\U1/aes_core/SB0/n518 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U219  ( .A(\U1/aes_core/SB0/n487 ), .B(
        \U1/aes_core/SB0/n524 ), .Y(\U1/aes_core/SB0/n520 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U218  ( .A(\U1/aes_core/SB0/n523 ), .B(
        \U1/aes_core/SB0/n482 ), .Y(\U1/aes_core/SB0/n521 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U217  ( .A0(\U1/aes_core/SB0/n520 ), 
        .A1(\U1/aes_core/SB0/n400 ), .B0(\U1/aes_core/SB0/n521 ), .B1(
        \U1/aes_core/SB0/n436 ), .C0(\U1/aes_core/SB0/n522 ), .C1(
        \U1/aes_core/SB0/n435 ), .Y(\U1/aes_core/SB0/n519 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U216  ( .A(\U1/aes_core/SB0/n427 ), .B(
        \U1/aes_core/SB0/n472 ), .C(\U1/aes_core/SB0/n516 ), .D(
        \U1/aes_core/SB0/n517 ), .E(\U1/aes_core/SB0/n518 ), .F(
        \U1/aes_core/SB0/n519 ), .Y(\U1/aes_core/sb0 [28]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U215  ( .A1N(\U1/aes_core/SB0/n514 ), 
        .A0(\U1/aes_core/SB0/n515 ), .B0(\U1/aes_core/SB0/n437 ), .Y(
        \U1/aes_core/SB0/n498 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U214  ( .A(\U1/aes_core/SB0/n424 ), .B(
        \U1/aes_core/SB0/n443 ), .Y(\U1/aes_core/SB0/n511 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U213  ( .A0(\U1/aes_core/SB0/n400 ), 
        .A1(\U1/aes_core/SB0/n510 ), .B0(\U1/aes_core/SB0/n511 ), .B1(
        \U1/aes_core/SB0/n397 ), .C0(\U1/aes_core/SB0/n512 ), .C1(
        \U1/aes_core/SB0/n513 ), .Y(\U1/aes_core/SB0/n499 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U212  ( .A(\U1/aes_core/SB0/n509 ), .Y(
        \U1/aes_core/SB0/n506 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U211  ( .AN(\U1/aes_core/SB0/n505 ), .B(
        \U1/aes_core/SB0/n506 ), .C(\U1/aes_core/SB0/n507 ), .D(
        \U1/aes_core/SB0/n508 ), .Y(\U1/aes_core/SB0/n500 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U210  ( .A(\U1/aes_core/SB0/n502 ), .B(
        \U1/aes_core/SB0/n503 ), .C(\U1/aes_core/SB0/n504 ), .Y(
        \U1/aes_core/SB0/n501 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U209  ( .A(\U1/aes_core/SB0/n496 ), .B(
        \U1/aes_core/SB0/n497 ), .C(\U1/aes_core/SB0/n498 ), .D(
        \U1/aes_core/SB0/n499 ), .E(\U1/aes_core/SB0/n500 ), .F(
        \U1/aes_core/SB0/n501 ), .Y(\U1/aes_core/SB0/n426 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U208  ( .A(\U1/aes_core/SB0/n495 ), .Y(
        \U1/aes_core/SB0/n493 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U207  ( .A0(\U1/aes_core/SB0/n413 ), .A1(
        \U1/aes_core/SB0/n416 ), .B0(\U1/aes_core/SB0/n412 ), .B1(
        \U1/aes_core/SB0/n414 ), .Y(\U1/aes_core/SB0/n494 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U206  ( .A0(\U1/aes_core/SB0/n437 ), 
        .A1(\U1/aes_core/SB0/n492 ), .B0(\U1/aes_core/SB0/n493 ), .C0(
        \U1/aes_core/SB0/n494 ), .Y(\U1/aes_core/SB0/n473 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U205  ( .A0(\U1/aes_core/SB0/n490 ), .A1(
        \U1/aes_core/SB0/n413 ), .B0(\U1/aes_core/SB0/n491 ), .Y(
        \U1/aes_core/SB0/n484 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U204  ( .A0(\U1/aes_core/SB0/n487 ), .A1(
        \U1/aes_core/SB0/n488 ), .B0(\U1/aes_core/SB0/n489 ), .Y(
        \U1/aes_core/SB0/n485 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U203  ( .AN(\U1/aes_core/SB0/n483 ), .B(
        \U1/aes_core/SB0/n484 ), .C(\U1/aes_core/SB0/n485 ), .D(
        \U1/aes_core/SB0/n486 ), .Y(\U1/aes_core/SB0/n474 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U202  ( .A0(\U1/aes_core/SB0/n417 ), .A1(
        \U1/aes_core/SB0/n481 ), .B0(\U1/aes_core/SB0/n482 ), .Y(
        \U1/aes_core/SB0/n477 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB0/U201  ( .A0(\U1/aes_core/SB0/n435 ), .A1(
        \U1/aes_core/SB0/n479 ), .B0(\U1/aes_core/SB0/n398 ), .B1(
        \U1/aes_core/SB0/n480 ), .Y(\U1/aes_core/SB0/n478 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U200  ( .A0(\U1/aes_core/SB0/n476 ), 
        .A1(\U1/aes_core/SB0/n436 ), .B0(\U1/aes_core/SB0/n477 ), .C0(
        \U1/aes_core/SB0/n478 ), .Y(\U1/aes_core/SB0/n475 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U199  ( .A(\U1/aes_core/SB0/n426 ), .B(
        \U1/aes_core/SB0/n471 ), .C(\U1/aes_core/SB0/n472 ), .D(
        \U1/aes_core/SB0/n473 ), .E(\U1/aes_core/SB0/n474 ), .F(
        \U1/aes_core/SB0/n475 ), .Y(\U1/aes_core/sb0 [29]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U198  ( .A0(\U1/aes_core/SB0/n142 ), .A1(
        \U1/aes_core/SB0/n122 ), .B0(\U1/aes_core/SB0/n101 ), .B1(
        \U1/aes_core/SB0/n111 ), .Y(\U1/aes_core/SB0/n470 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U197  ( .A0(\U1/aes_core/SB0/n191 ), 
        .A1(\U1/aes_core/SB0/n97 ), .B0(\U1/aes_core/SB0/n241 ), .B1(
        \U1/aes_core/SB0/n170 ), .C0(\U1/aes_core/SB0/n470 ), .Y(
        \U1/aes_core/SB0/n464 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U196  ( .A(\U1/aes_core/SB0/n116 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n307 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U195  ( .A(\U1/aes_core/SB0/n142 ), .B(
        \U1/aes_core/SB0/n166 ), .Y(\U1/aes_core/SB0/n326 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U194  ( .A(\U1/aes_core/SB0/n122 ), .B(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n358 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U193  ( .A(\U1/aes_core/SB0/n202 ), .B(
        \U1/aes_core/SB0/n159 ), .Y(\U1/aes_core/SB0/n339 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U192  ( .A(\U1/aes_core/SB0/n307 ), .B(
        \U1/aes_core/SB0/n326 ), .C(\U1/aes_core/SB0/n358 ), .D(
        \U1/aes_core/SB0/n339 ), .Y(\U1/aes_core/SB0/n465 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U191  ( .A(\U1/aes_core/SB0/n96 ), .B(
        \U1/aes_core/SB0/n118 ), .Y(\U1/aes_core/SB0/n213 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U190  ( .A0(\U1/aes_core/SB0/n165 ), .A1(
        \U1/aes_core/SB0/n213 ), .B0(\U1/aes_core/SB0/n112 ), .Y(
        \U1/aes_core/SB0/n467 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U189  ( .A0(\U1/aes_core/SB0/n115 ), .A1(
        \U1/aes_core/SB0/n224 ), .B0(\U1/aes_core/SB0/n212 ), .Y(
        \U1/aes_core/SB0/n468 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U188  ( .A0(\U1/aes_core/SB0/n207 ), .A1(
        \U1/aes_core/SB0/n167 ), .B0(\U1/aes_core/SB0/n113 ), .Y(
        \U1/aes_core/SB0/n469 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U187  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n115 ), .Y(\U1/aes_core/SB0/n240 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U186  ( .A(\U1/aes_core/SB0/n467 ), .B(
        \U1/aes_core/SB0/n468 ), .C(\U1/aes_core/SB0/n469 ), .D(
        \U1/aes_core/SB0/n240 ), .Y(\U1/aes_core/SB0/n466 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U185  ( .A(\U1/aes_core/SB0/n461 ), .B(
        \U1/aes_core/SB0/n462 ), .C(\U1/aes_core/SB0/n463 ), .D(
        \U1/aes_core/SB0/n464 ), .E(\U1/aes_core/SB0/n465 ), .F(
        \U1/aes_core/SB0/n466 ), .Y(\U1/aes_core/SB0/n92 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U184  ( .A0(\U1/aes_core/SB0/n286 ), 
        .A1(\U1/aes_core/SB0/n111 ), .B0(\U1/aes_core/SB0/n103 ), .B1(
        \U1/aes_core/SB0/n168 ), .C0(\U1/aes_core/SB0/n92 ), .Y(
        \U1/aes_core/SB0/n460 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U183  ( .A(\U1/aes_core/SB0/n460 ), .Y(
        \U1/aes_core/SB0/n453 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U182  ( .A(\U1/aes_core/SB0/n159 ), .B(
        \U1/aes_core/SB0/n372 ), .Y(\U1/aes_core/SB0/n250 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U181  ( .A1N(\U1/aes_core/SB0/n250 ), 
        .A0(\U1/aes_core/SB0/n141 ), .B0(\U1/aes_core/SB0/n169 ), .Y(
        \U1/aes_core/SB0/n457 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U180  ( .A0(\U1/aes_core/SB0/n201 ), .A1(
        \U1/aes_core/SB0/n293 ), .B0(\U1/aes_core/SB0/n142 ), .Y(
        \U1/aes_core/SB0/n458 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U179  ( .A0(\U1/aes_core/SB0/n115 ), .A1(
        \U1/aes_core/SB0/n160 ), .B0(\U1/aes_core/SB0/n121 ), .Y(
        \U1/aes_core/SB0/n459 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U178  ( .A(\U1/aes_core/SB0/n144 ), .B(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n343 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U177  ( .A(\U1/aes_core/SB0/n457 ), .B(
        \U1/aes_core/SB0/n458 ), .C(\U1/aes_core/SB0/n459 ), .D(
        \U1/aes_core/SB0/n343 ), .Y(\U1/aes_core/SB0/n454 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U176  ( .A(\U1/aes_core/SB0/n145 ), .B(
        \U1/aes_core/SB0/n113 ), .Y(\U1/aes_core/SB0/n114 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U175  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n167 ), .Y(\U1/aes_core/SB0/n456 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U174  ( .A0(\U1/aes_core/SB0/n114 ), 
        .A1(\U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n456 ), .B1(
        \U1/aes_core/SB0/n133 ), .C0(\U1/aes_core/SB0/n190 ), .C1(
        \U1/aes_core/SB0/n188 ), .Y(\U1/aes_core/SB0/n455 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U173  ( .A(\U1/aes_core/SB0/n450 ), .B(
        \U1/aes_core/SB0/n451 ), .C(\U1/aes_core/SB0/n452 ), .D(
        \U1/aes_core/SB0/n453 ), .E(\U1/aes_core/SB0/n454 ), .F(
        \U1/aes_core/SB0/n455 ), .Y(\U1/aes_core/sb0 [2]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U172  ( .A0(\U1/aes_core/SB0/n447 ), 
        .A1(\U1/aes_core/SB0/n407 ), .B0(\U1/aes_core/SB0/n448 ), .B1(
        \U1/aes_core/SB0/n400 ), .C0(\U1/aes_core/SB0/n449 ), .Y(
        \U1/aes_core/SB0/n429 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U171  ( .A0(\U1/aes_core/SB0/n446 ), .A1(
        \U1/aes_core/SB0/n402 ), .B0(\U1/aes_core/SB0/n413 ), .Y(
        \U1/aes_core/SB0/n438 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U170  ( .A0(\U1/aes_core/SB0/n422 ), .A1(
        \U1/aes_core/SB0/n445 ), .B0(\U1/aes_core/SB0/n414 ), .Y(
        \U1/aes_core/SB0/n439 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U169  ( .A0(\U1/aes_core/SB0/n442 ), .A1(
        \U1/aes_core/SB0/n443 ), .B0(\U1/aes_core/SB0/n444 ), .Y(
        \U1/aes_core/SB0/n440 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U168  ( .A(\U1/aes_core/SB0/n438 ), .B(
        \U1/aes_core/SB0/n439 ), .C(\U1/aes_core/SB0/n440 ), .D(
        \U1/aes_core/SB0/n441 ), .Y(\U1/aes_core/SB0/n430 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U167  ( .A(\U1/aes_core/SB0/n407 ), .B(
        \U1/aes_core/SB0/n437 ), .Y(\U1/aes_core/SB0/n405 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U166  ( .A(\U1/aes_core/SB0/n417 ), .B(
        \U1/aes_core/SB0/n405 ), .Y(\U1/aes_core/SB0/n433 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U165  ( .A0(\U1/aes_core/SB0/n419 ), 
        .A1(\U1/aes_core/SB0/n432 ), .B0(\U1/aes_core/SB0/n433 ), .B1(
        \U1/aes_core/SB0/n434 ), .C0(\U1/aes_core/SB0/n435 ), .C1(
        \U1/aes_core/SB0/n436 ), .Y(\U1/aes_core/SB0/n431 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U164  ( .A(\U1/aes_core/SB0/n426 ), .B(
        \U1/aes_core/SB0/n427 ), .C(\U1/aes_core/SB0/n428 ), .D(
        \U1/aes_core/SB0/n429 ), .E(\U1/aes_core/SB0/n430 ), .F(
        \U1/aes_core/SB0/n431 ), .Y(\U1/aes_core/sb0 [30]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U163  ( .A0(\U1/aes_core/SB0/n422 ), .A1(
        \U1/aes_core/SB0/n423 ), .B0(\U1/aes_core/SB0/n424 ), .B1(
        \U1/aes_core/SB0/n425 ), .Y(\U1/aes_core/SB0/n421 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U162  ( .A0(\U1/aes_core/SB0/n418 ), 
        .A1(\U1/aes_core/SB0/n419 ), .B0(\U1/aes_core/SB0/n420 ), .C0(
        \U1/aes_core/SB0/n421 ), .Y(\U1/aes_core/SB0/n394 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U161  ( .A1N(\U1/aes_core/SB0/n415 ), 
        .A0(\U1/aes_core/SB0/n416 ), .B0(\U1/aes_core/SB0/n417 ), .Y(
        \U1/aes_core/SB0/n408 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U160  ( .A0(\U1/aes_core/SB0/n412 ), .A1(
        \U1/aes_core/SB0/n413 ), .B0(\U1/aes_core/SB0/n414 ), .Y(
        \U1/aes_core/SB0/n409 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U159  ( .A(\U1/aes_core/SB0/n408 ), .B(
        \U1/aes_core/SB0/n409 ), .C(\U1/aes_core/SB0/n410 ), .D(
        \U1/aes_core/SB0/n411 ), .Y(\U1/aes_core/SB0/n395 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U158  ( .A(\U1/aes_core/SB0/n406 ), .B(
        \U1/aes_core/SB0/n407 ), .Y(\U1/aes_core/SB0/n403 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U157  ( .A0(\U1/aes_core/SB0/n402 ), .A1(
        \U1/aes_core/SB0/n403 ), .B0(\U1/aes_core/SB0/n404 ), .B1(
        \U1/aes_core/SB0/n405 ), .Y(\U1/aes_core/SB0/n401 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U156  ( .A0(\U1/aes_core/SB0/n397 ), 
        .A1(\U1/aes_core/SB0/n398 ), .B0(\U1/aes_core/SB0/n399 ), .B1(
        \U1/aes_core/SB0/n400 ), .C0(\U1/aes_core/SB0/n401 ), .Y(
        \U1/aes_core/SB0/n396 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U155  ( .A(\U1/aes_core/SB0/n391 ), .B(
        \U1/aes_core/SB0/n392 ), .C(\U1/aes_core/SB0/n393 ), .D(
        \U1/aes_core/SB0/n394 ), .E(\U1/aes_core/SB0/n395 ), .F(
        \U1/aes_core/SB0/n396 ), .Y(\U1/aes_core/sb0 [31]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U154  ( .A(\U1/aes_core/SB0/n286 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n109 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U153  ( .AN(\U1/aes_core/SB0/n388 ), .B(
        \U1/aes_core/SB0/n389 ), .C(\U1/aes_core/SB0/n390 ), .D(
        \U1/aes_core/SB0/n109 ), .Y(\U1/aes_core/SB0/n380 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U152  ( .A0(\U1/aes_core/SB0/n387 ), .A1(
        \U1/aes_core/SB0/n142 ), .B0(\U1/aes_core/SB0/n224 ), .Y(
        \U1/aes_core/SB0/n384 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U149  ( .A(\U1/aes_core/SB0/n168 ), .B(
        \U1/aes_core/SB0/n121 ), .Y(\U1/aes_core/SB0/n157 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U148  ( .A0(\U1/aes_core/SB0/n278 ), 
        .A1(\U1/aes_core/SB0/n99 ), .B0(\U1/aes_core/SB0/n157 ), .B1(
        \U1/aes_core/SB0/n146 ), .C0(\U1/aes_core/SB0/n105 ), .C1(
        \U1/aes_core/SB0/n96 ), .Y(\U1/aes_core/SB0/n382 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U147  ( .A(\U1/aes_core/SB0/n377 ), .B(
        \U1/aes_core/SB0/n378 ), .C(\U1/aes_core/SB0/n379 ), .D(
        \U1/aes_core/SB0/n380 ), .E(\U1/aes_core/SB0/n381 ), .F(
        \U1/aes_core/SB0/n382 ), .Y(\U1/aes_core/SB0/n194 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U146  ( .AN(\U1/aes_core/SB0/n373 ), .B(
        \U1/aes_core/SB0/n374 ), .C(\U1/aes_core/SB0/n375 ), .D(
        \U1/aes_core/SB0/n376 ), .Y(\U1/aes_core/SB0/n363 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB0/U145  ( .A0(\U1/aes_core/SB0/n111 ), 
        .A1(\U1/aes_core/SB0/n201 ), .B0(\U1/aes_core/SB0/n116 ), .B1(
        \U1/aes_core/SB0/n202 ), .C0(\U1/aes_core/SB0/n372 ), .C1(
        \U1/aes_core/SB0/n101 ), .Y(\U1/aes_core/SB0/n364 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U144  ( .A0(\U1/aes_core/SB0/n147 ), .A1(
        \U1/aes_core/SB0/n241 ), .B0(\U1/aes_core/SB0/n371 ), .B1(
        \U1/aes_core/SB0/n278 ), .Y(\U1/aes_core/SB0/n370 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U143  ( .A0(\U1/aes_core/SB0/n224 ), 
        .A1(\U1/aes_core/SB0/n207 ), .B0(\U1/aes_core/SB0/n208 ), .B1(
        \U1/aes_core/SB0/n144 ), .C0(\U1/aes_core/SB0/n370 ), .Y(
        \U1/aes_core/SB0/n365 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U142  ( .A(\U1/aes_core/SB0/n136 ), .B(
        \U1/aes_core/SB0/n97 ), .Y(\U1/aes_core/SB0/n368 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U141  ( .A0(\U1/aes_core/SB0/n286 ), 
        .A1(\U1/aes_core/SB0/n367 ), .B0(\U1/aes_core/SB0/n115 ), .B1(
        \U1/aes_core/SB0/n368 ), .C0(\U1/aes_core/SB0/n369 ), .Y(
        \U1/aes_core/SB0/n366 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U140  ( .AN(\U1/aes_core/SB0/n363 ), .B(
        \U1/aes_core/SB0/n364 ), .C(\U1/aes_core/SB0/n365 ), .D(
        \U1/aes_core/SB0/n366 ), .Y(\U1/aes_core/SB0/n149 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U139  ( .A(\U1/aes_core/SB0/n362 ), .Y(
        \U1/aes_core/SB0/n346 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U138  ( .A0(\U1/aes_core/SB0/n257 ), .A1(
        \U1/aes_core/SB0/n188 ), .B0(\U1/aes_core/SB0/n361 ), .Y(
        \U1/aes_core/SB0/n347 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U137  ( .A0(\U1/aes_core/SB0/n115 ), .A1(
        \U1/aes_core/SB0/n116 ), .B0(\U1/aes_core/SB0/n145 ), .B1(
        \U1/aes_core/SB0/n360 ), .Y(\U1/aes_core/SB0/n359 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U136  ( .A0(\U1/aes_core/SB0/n134 ), 
        .A1(\U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n118 ), .B1(
        \U1/aes_core/SB0/n106 ), .C0(\U1/aes_core/SB0/n359 ), .Y(
        \U1/aes_core/SB0/n348 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U135  ( .A(\U1/aes_core/SB0/n355 ), .B(
        \U1/aes_core/SB0/n356 ), .C(\U1/aes_core/SB0/n357 ), .D(
        \U1/aes_core/SB0/n358 ), .Y(\U1/aes_core/SB0/n349 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U134  ( .AN(\U1/aes_core/SB0/n351 ), .B(
        \U1/aes_core/SB0/n352 ), .C(\U1/aes_core/SB0/n353 ), .D(
        \U1/aes_core/SB0/n354 ), .Y(\U1/aes_core/SB0/n350 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U133  ( .A(\U1/aes_core/SB0/n345 ), .B(
        \U1/aes_core/SB0/n346 ), .C(\U1/aes_core/SB0/n347 ), .D(
        \U1/aes_core/SB0/n348 ), .E(\U1/aes_core/SB0/n349 ), .F(
        \U1/aes_core/SB0/n350 ), .Y(\U1/aes_core/SB0/n245 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U132  ( .A0(\U1/aes_core/SB0/n158 ), .A1(
        \U1/aes_core/SB0/n241 ), .B0(\U1/aes_core/SB0/n344 ), .Y(
        \U1/aes_core/SB0/n329 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U131  ( .AN(\U1/aes_core/SB0/n340 ), .B(
        \U1/aes_core/SB0/n341 ), .C(\U1/aes_core/SB0/n342 ), .D(
        \U1/aes_core/SB0/n343 ), .Y(\U1/aes_core/SB0/n330 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U130  ( .A(\U1/aes_core/SB0/n124 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n110 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U129  ( .A(\U1/aes_core/SB0/n337 ), .B(
        \U1/aes_core/SB0/n338 ), .C(\U1/aes_core/SB0/n339 ), .D(
        \U1/aes_core/SB0/n110 ), .Y(\U1/aes_core/SB0/n331 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U128  ( .A(\U1/aes_core/SB0/n333 ), .B(
        \U1/aes_core/SB0/n334 ), .C(\U1/aes_core/SB0/n335 ), .D(
        \U1/aes_core/SB0/n336 ), .Y(\U1/aes_core/SB0/n332 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U127  ( .A(\U1/aes_core/SB0/n327 ), .B(
        \U1/aes_core/SB0/n328 ), .C(\U1/aes_core/SB0/n329 ), .D(
        \U1/aes_core/SB0/n330 ), .E(\U1/aes_core/SB0/n331 ), .F(
        \U1/aes_core/SB0/n332 ), .Y(\U1/aes_core/SB0/n221 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U126  ( .AN(\U1/aes_core/SB0/n323 ), .B(
        \U1/aes_core/SB0/n324 ), .C(\U1/aes_core/SB0/n325 ), .D(
        \U1/aes_core/SB0/n326 ), .Y(\U1/aes_core/SB0/n314 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U125  ( .A(\U1/aes_core/SB0/n319 ), .B(
        \U1/aes_core/SB0/n320 ), .C(\U1/aes_core/SB0/n321 ), .D(
        \U1/aes_core/SB0/n322 ), .Y(\U1/aes_core/SB0/n315 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U124  ( .A(\U1/aes_core/SB0/n159 ), .B(
        \U1/aes_core/SB0/n123 ), .C(\U1/aes_core/SB0/n121 ), .Y(
        \U1/aes_core/SB0/n317 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U123  ( .A0(\U1/aes_core/SB0/n317 ), 
        .A1(\U1/aes_core/SB0/n133 ), .B0(\U1/aes_core/SB0/n278 ), .B1(
        \U1/aes_core/SB0/n97 ), .C0(\U1/aes_core/SB0/n318 ), .Y(
        \U1/aes_core/SB0/n316 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U122  ( .A(\U1/aes_core/SB0/n311 ), .B(
        \U1/aes_core/SB0/n312 ), .C(\U1/aes_core/SB0/n313 ), .D(
        \U1/aes_core/SB0/n314 ), .E(\U1/aes_core/SB0/n315 ), .F(
        \U1/aes_core/SB0/n316 ), .Y(\U1/aes_core/SB0/n173 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U121  ( .A0(\U1/aes_core/SB0/n278 ), .A1(
        \U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n310 ), .Y(
        \U1/aes_core/SB0/n296 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U120  ( .A0(\U1/aes_core/SB0/n169 ), .A1(
        \U1/aes_core/SB0/n167 ), .B0(\U1/aes_core/SB0/n112 ), .B1(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n309 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U119  ( .A0(\U1/aes_core/SB0/n258 ), 
        .A1(\U1/aes_core/SB0/n170 ), .B0(\U1/aes_core/SB0/n257 ), .B1(
        \U1/aes_core/SB0/n193 ), .C0(\U1/aes_core/SB0/n309 ), .Y(
        \U1/aes_core/SB0/n297 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U118  ( .A(\U1/aes_core/SB0/n308 ), .Y(
        \U1/aes_core/SB0/n305 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U117  ( .AN(\U1/aes_core/SB0/n304 ), .B(
        \U1/aes_core/SB0/n305 ), .C(\U1/aes_core/SB0/n306 ), .D(
        \U1/aes_core/SB0/n307 ), .Y(\U1/aes_core/SB0/n298 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U116  ( .A(\U1/aes_core/SB0/n300 ), .B(
        \U1/aes_core/SB0/n301 ), .C(\U1/aes_core/SB0/n302 ), .D(
        \U1/aes_core/SB0/n303 ), .Y(\U1/aes_core/SB0/n299 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U115  ( .A(\U1/aes_core/SB0/n294 ), .B(
        \U1/aes_core/SB0/n295 ), .C(\U1/aes_core/SB0/n296 ), .D(
        \U1/aes_core/SB0/n297 ), .E(\U1/aes_core/SB0/n298 ), .F(
        \U1/aes_core/SB0/n299 ), .Y(\U1/aes_core/SB0/n214 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U114  ( .A0(\U1/aes_core/SB0/n123 ), .A1(
        \U1/aes_core/SB0/n293 ), .B0(\U1/aes_core/SB0/n113 ), .B1(
        \U1/aes_core/SB0/n167 ), .Y(\U1/aes_core/SB0/n292 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U113  ( .A0(\U1/aes_core/SB0/n241 ), 
        .A1(\U1/aes_core/SB0/n96 ), .B0(\U1/aes_core/SB0/n291 ), .B1(
        \U1/aes_core/SB0/n106 ), .C0(\U1/aes_core/SB0/n292 ), .Y(
        \U1/aes_core/SB0/n279 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U112  ( .AN(\U1/aes_core/SB0/n287 ), .B(
        \U1/aes_core/SB0/n288 ), .C(\U1/aes_core/SB0/n289 ), .D(
        \U1/aes_core/SB0/n290 ), .Y(\U1/aes_core/SB0/n280 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U111  ( .A0(\U1/aes_core/SB0/n103 ), .A1(
        \U1/aes_core/SB0/n286 ), .B0(\U1/aes_core/SB0/n112 ), .Y(
        \U1/aes_core/SB0/n282 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U110  ( .A(\U1/aes_core/SB0/n136 ), .B(
        \U1/aes_core/SB0/n131 ), .Y(\U1/aes_core/SB0/n285 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U109  ( .A0(\U1/aes_core/SB0/n160 ), .A1(
        \U1/aes_core/SB0/n285 ), .B0(\U1/aes_core/SB0/n159 ), .B1(
        \U1/aes_core/SB0/n213 ), .Y(\U1/aes_core/SB0/n284 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U108  ( .A(\U1/aes_core/SB0/n282 ), .B(
        \U1/aes_core/SB0/n283 ), .C(\U1/aes_core/SB0/n284 ), .Y(
        \U1/aes_core/SB0/n281 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U107  ( .A(\U1/aes_core/SB0/n221 ), .B(
        \U1/aes_core/SB0/n173 ), .C(\U1/aes_core/SB0/n214 ), .D(
        \U1/aes_core/SB0/n279 ), .E(\U1/aes_core/SB0/n280 ), .F(
        \U1/aes_core/SB0/n281 ), .Y(\U1/aes_core/SB0/n127 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U106  ( .A(\U1/aes_core/SB0/n194 ), .B(
        \U1/aes_core/SB0/n149 ), .C(\U1/aes_core/SB0/n245 ), .D(
        \U1/aes_core/SB0/n127 ), .Y(\U1/aes_core/SB0/n265 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U105  ( .A0(\U1/aes_core/SB0/n147 ), .A1(
        \U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n278 ), .B1(
        \U1/aes_core/SB0/n131 ), .Y(\U1/aes_core/SB0/n277 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U104  ( .A0(\U1/aes_core/SB0/n142 ), 
        .A1(\U1/aes_core/SB0/n124 ), .B0(\U1/aes_core/SB0/n111 ), .B1(
        \U1/aes_core/SB0/n103 ), .C0(\U1/aes_core/SB0/n277 ), .Y(
        \U1/aes_core/SB0/n266 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U103  ( .A(\U1/aes_core/SB0/n276 ), .Y(
        \U1/aes_core/SB0/n273 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U102  ( .A0(\U1/aes_core/SB0/n275 ), .A1(
        \U1/aes_core/SB0/n170 ), .B0(\U1/aes_core/SB0/n242 ), .B1(
        \U1/aes_core/SB0/n190 ), .Y(\U1/aes_core/SB0/n274 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U101  ( .A0(\U1/aes_core/SB0/n123 ), 
        .A1(\U1/aes_core/SB0/n273 ), .B0(\U1/aes_core/SB0/n141 ), .B1(
        \U1/aes_core/SB0/n192 ), .C0(\U1/aes_core/SB0/n274 ), .Y(
        \U1/aes_core/SB0/n267 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U100  ( .A0(\U1/aes_core/SB0/n101 ), .A1(
        \U1/aes_core/SB0/n224 ), .B0(\U1/aes_core/SB0/n121 ), .Y(
        \U1/aes_core/SB0/n269 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB0/U99  ( .A(\U1/aes_core/SB0/n269 ), .B(
        \U1/aes_core/SB0/n270 ), .C(\U1/aes_core/SB0/n271 ), .D(
        \U1/aes_core/SB0/n272 ), .Y(\U1/aes_core/SB0/n268 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U98  ( .AN(\U1/aes_core/SB0/n265 ), .B(
        \U1/aes_core/SB0/n266 ), .C(\U1/aes_core/SB0/n267 ), .D(
        \U1/aes_core/SB0/n268 ), .Y(\U1/aes_core/sb0 [3]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U97  ( .A0(\U1/aes_core/SB0/n250 ), .A1(
        \U1/aes_core/SB0/n135 ), .B0(\U1/aes_core/SB0/n191 ), .Y(
        \U1/aes_core/SB0/n253 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U96  ( .A(\U1/aes_core/SB0/n262 ), .B(
        \U1/aes_core/SB0/n263 ), .C(\U1/aes_core/SB0/n264 ), .Y(
        \U1/aes_core/SB0/n254 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U95  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n112 ), .Y(\U1/aes_core/SB0/n259 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U94  ( .A(\U1/aes_core/SB0/n141 ), .B(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n261 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U93  ( .A0(\U1/aes_core/SB0/n259 ), .A1(
        \U1/aes_core/SB0/n260 ), .B0(\U1/aes_core/SB0/n261 ), .B1(
        \U1/aes_core/SB0/n118 ), .C0(\U1/aes_core/SB0/n135 ), .C1(
        \U1/aes_core/SB0/n209 ), .Y(\U1/aes_core/SB0/n255 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U92  ( .A0(\U1/aes_core/SB0/n158 ), .A1(
        \U1/aes_core/SB0/n257 ), .B0(\U1/aes_core/SB0/n96 ), .B1(
        \U1/aes_core/SB0/n106 ), .C0(\U1/aes_core/SB0/n133 ), .C1(
        \U1/aes_core/SB0/n258 ), .Y(\U1/aes_core/SB0/n256 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U91  ( .A(\U1/aes_core/SB0/n251 ), .B(
        \U1/aes_core/SB0/n252 ), .C(\U1/aes_core/SB0/n253 ), .D(
        \U1/aes_core/SB0/n254 ), .E(\U1/aes_core/SB0/n255 ), .F(
        \U1/aes_core/SB0/n256 ), .Y(\U1/aes_core/SB0/n126 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB0/U90  ( .A0(\U1/aes_core/SB0/n250 ), .A1(
        \U1/aes_core/SB0/n241 ), .B0(\U1/aes_core/SB0/n170 ), .Y(
        \U1/aes_core/SB0/n215 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB0/U89  ( .A0(\U1/aes_core/SB0/n146 ), .A1(
        \U1/aes_core/SB0/n133 ), .A2(\U1/aes_core/SB0/n193 ), .B0(
        \U1/aes_core/SB0/n117 ), .Y(\U1/aes_core/SB0/n216 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U88  ( .A(\U1/aes_core/SB0/n246 ), .B(
        \U1/aes_core/SB0/n247 ), .C(\U1/aes_core/SB0/n248 ), .D(
        \U1/aes_core/SB0/n249 ), .Y(\U1/aes_core/SB0/n219 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U87  ( .A(\U1/aes_core/SB0/n245 ), .Y(
        \U1/aes_core/SB0/n222 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U86  ( .A(\U1/aes_core/SB0/n244 ), .Y(
        \U1/aes_core/SB0/n228 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB0/U85  ( .A0(\U1/aes_core/SB0/n242 ), .A1(
        \U1/aes_core/SB0/n105 ), .B0N(\U1/aes_core/SB0/n243 ), .Y(
        \U1/aes_core/SB0/n229 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U84  ( .A0(\U1/aes_core/SB0/n98 ), .A1(
        \U1/aes_core/SB0/n241 ), .B0(\U1/aes_core/SB0/n191 ), .B1(
        \U1/aes_core/SB0/n131 ), .C0(\U1/aes_core/SB0/n117 ), .C1(
        \U1/aes_core/SB0/n96 ), .Y(\U1/aes_core/SB0/n230 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U83  ( .AN(\U1/aes_core/SB0/n237 ), .B(
        \U1/aes_core/SB0/n238 ), .C(\U1/aes_core/SB0/n239 ), .D(
        \U1/aes_core/SB0/n240 ), .Y(\U1/aes_core/SB0/n231 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U82  ( .A(\U1/aes_core/SB0/n233 ), .B(
        \U1/aes_core/SB0/n234 ), .C(\U1/aes_core/SB0/n235 ), .D(
        \U1/aes_core/SB0/n236 ), .Y(\U1/aes_core/SB0/n232 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U81  ( .A(\U1/aes_core/SB0/n227 ), .B(
        \U1/aes_core/SB0/n228 ), .C(\U1/aes_core/SB0/n229 ), .D(
        \U1/aes_core/SB0/n230 ), .E(\U1/aes_core/SB0/n231 ), .F(
        \U1/aes_core/SB0/n232 ), .Y(\U1/aes_core/SB0/n226 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U80  ( .A(\U1/aes_core/SB0/n226 ), .Y(
        \U1/aes_core/SB0/n148 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U79  ( .A0(\U1/aes_core/SB0/n158 ), .A1(
        \U1/aes_core/SB0/n136 ), .B0(\U1/aes_core/SB0/n96 ), .B1(
        \U1/aes_core/SB0/n97 ), .Y(\U1/aes_core/SB0/n225 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U78  ( .A0(\U1/aes_core/SB0/n168 ), .A1(
        \U1/aes_core/SB0/n224 ), .B0(\U1/aes_core/SB0/n144 ), .B1(
        \U1/aes_core/SB0/n122 ), .C0(\U1/aes_core/SB0/n225 ), .Y(
        \U1/aes_core/SB0/n223 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U77  ( .AN(\U1/aes_core/SB0/n221 ), .B(
        \U1/aes_core/SB0/n222 ), .C(\U1/aes_core/SB0/n148 ), .D(
        \U1/aes_core/SB0/n223 ), .Y(\U1/aes_core/SB0/n220 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U76  ( .A(\U1/aes_core/SB0/n215 ), .B(
        \U1/aes_core/SB0/n216 ), .C(\U1/aes_core/SB0/n217 ), .D(
        \U1/aes_core/SB0/n218 ), .E(\U1/aes_core/SB0/n219 ), .F(
        \U1/aes_core/SB0/n220 ), .Y(\U1/aes_core/SB0/n150 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U75  ( .A(\U1/aes_core/SB0/n214 ), .Y(
        \U1/aes_core/SB0/n210 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U74  ( .A0(\U1/aes_core/SB0/n212 ), .A1(
        \U1/aes_core/SB0/n213 ), .B0(\U1/aes_core/SB0/n166 ), .B1(
        \U1/aes_core/SB0/n207 ), .Y(\U1/aes_core/SB0/n211 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U73  ( .A0(\U1/aes_core/SB0/n117 ), .A1(
        \U1/aes_core/SB0/n209 ), .B0(\U1/aes_core/SB0/n210 ), .C0(
        \U1/aes_core/SB0/n211 ), .Y(\U1/aes_core/SB0/n195 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U72  ( .A0(\U1/aes_core/SB0/n208 ), .A1(
        \U1/aes_core/SB0/n145 ), .B0(\U1/aes_core/SB0/n116 ), .Y(
        \U1/aes_core/SB0/n203 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U71  ( .A0(\U1/aes_core/SB0/n207 ), .A1(
        \U1/aes_core/SB0/n142 ), .B0(\U1/aes_core/SB0/n113 ), .Y(
        \U1/aes_core/SB0/n204 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U70  ( .A(\U1/aes_core/SB0/n203 ), .B(
        \U1/aes_core/SB0/n204 ), .C(\U1/aes_core/SB0/n205 ), .D(
        \U1/aes_core/SB0/n206 ), .Y(\U1/aes_core/SB0/n196 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U69  ( .A(\U1/aes_core/SB0/n165 ), .B(
        \U1/aes_core/SB0/n202 ), .Y(\U1/aes_core/SB0/n198 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U68  ( .A(\U1/aes_core/SB0/n201 ), .B(
        \U1/aes_core/SB0/n160 ), .Y(\U1/aes_core/SB0/n199 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U67  ( .A0(\U1/aes_core/SB0/n198 ), .A1(
        \U1/aes_core/SB0/n99 ), .B0(\U1/aes_core/SB0/n199 ), .B1(
        \U1/aes_core/SB0/n135 ), .C0(\U1/aes_core/SB0/n200 ), .C1(
        \U1/aes_core/SB0/n134 ), .Y(\U1/aes_core/SB0/n197 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U66  ( .A(\U1/aes_core/SB0/n126 ), .B(
        \U1/aes_core/SB0/n150 ), .C(\U1/aes_core/SB0/n194 ), .D(
        \U1/aes_core/SB0/n195 ), .E(\U1/aes_core/SB0/n196 ), .F(
        \U1/aes_core/SB0/n197 ), .Y(\U1/aes_core/sb0 [4]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U65  ( .A1N(\U1/aes_core/SB0/n192 ), 
        .A0(\U1/aes_core/SB0/n193 ), .B0(\U1/aes_core/SB0/n136 ), .Y(
        \U1/aes_core/SB0/n176 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U64  ( .A(\U1/aes_core/SB0/n123 ), .B(
        \U1/aes_core/SB0/n142 ), .Y(\U1/aes_core/SB0/n189 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U63  ( .A0(\U1/aes_core/SB0/n99 ), .A1(
        \U1/aes_core/SB0/n188 ), .B0(\U1/aes_core/SB0/n189 ), .B1(
        \U1/aes_core/SB0/n96 ), .C0(\U1/aes_core/SB0/n190 ), .C1(
        \U1/aes_core/SB0/n191 ), .Y(\U1/aes_core/SB0/n177 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U62  ( .A(\U1/aes_core/SB0/n187 ), .Y(
        \U1/aes_core/SB0/n184 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U61  ( .AN(\U1/aes_core/SB0/n183 ), .B(
        \U1/aes_core/SB0/n184 ), .C(\U1/aes_core/SB0/n185 ), .D(
        \U1/aes_core/SB0/n186 ), .Y(\U1/aes_core/SB0/n178 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U60  ( .A(\U1/aes_core/SB0/n180 ), .B(
        \U1/aes_core/SB0/n181 ), .C(\U1/aes_core/SB0/n182 ), .Y(
        \U1/aes_core/SB0/n179 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U59  ( .A(\U1/aes_core/SB0/n174 ), .B(
        \U1/aes_core/SB0/n175 ), .C(\U1/aes_core/SB0/n176 ), .D(
        \U1/aes_core/SB0/n177 ), .E(\U1/aes_core/SB0/n178 ), .F(
        \U1/aes_core/SB0/n179 ), .Y(\U1/aes_core/SB0/n125 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U58  ( .A(\U1/aes_core/SB0/n173 ), .Y(
        \U1/aes_core/SB0/n171 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U57  ( .A0(\U1/aes_core/SB0/n112 ), .A1(
        \U1/aes_core/SB0/n115 ), .B0(\U1/aes_core/SB0/n111 ), .B1(
        \U1/aes_core/SB0/n113 ), .Y(\U1/aes_core/SB0/n172 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U56  ( .A0(\U1/aes_core/SB0/n136 ), .A1(
        \U1/aes_core/SB0/n170 ), .B0(\U1/aes_core/SB0/n171 ), .C0(
        \U1/aes_core/SB0/n172 ), .Y(\U1/aes_core/SB0/n151 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U55  ( .A0(\U1/aes_core/SB0/n168 ), .A1(
        \U1/aes_core/SB0/n112 ), .B0(\U1/aes_core/SB0/n169 ), .Y(
        \U1/aes_core/SB0/n162 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U54  ( .A0(\U1/aes_core/SB0/n165 ), .A1(
        \U1/aes_core/SB0/n166 ), .B0(\U1/aes_core/SB0/n167 ), .Y(
        \U1/aes_core/SB0/n163 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U53  ( .AN(\U1/aes_core/SB0/n161 ), .B(
        \U1/aes_core/SB0/n162 ), .C(\U1/aes_core/SB0/n163 ), .D(
        \U1/aes_core/SB0/n164 ), .Y(\U1/aes_core/SB0/n152 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U52  ( .A0(\U1/aes_core/SB0/n116 ), .A1(
        \U1/aes_core/SB0/n159 ), .B0(\U1/aes_core/SB0/n160 ), .Y(
        \U1/aes_core/SB0/n155 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB0/U51  ( .A0(\U1/aes_core/SB0/n134 ), .A1(
        \U1/aes_core/SB0/n157 ), .B0(\U1/aes_core/SB0/n97 ), .B1(
        \U1/aes_core/SB0/n158 ), .Y(\U1/aes_core/SB0/n156 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U50  ( .A0(\U1/aes_core/SB0/n154 ), .A1(
        \U1/aes_core/SB0/n135 ), .B0(\U1/aes_core/SB0/n155 ), .C0(
        \U1/aes_core/SB0/n156 ), .Y(\U1/aes_core/SB0/n153 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U49  ( .A(\U1/aes_core/SB0/n125 ), .B(
        \U1/aes_core/SB0/n149 ), .C(\U1/aes_core/SB0/n150 ), .D(
        \U1/aes_core/SB0/n151 ), .E(\U1/aes_core/SB0/n152 ), .F(
        \U1/aes_core/SB0/n153 ), .Y(\U1/aes_core/sb0 [5]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U48  ( .A0(\U1/aes_core/SB0/n146 ), .A1(
        \U1/aes_core/SB0/n106 ), .B0(\U1/aes_core/SB0/n147 ), .B1(
        \U1/aes_core/SB0/n99 ), .C0(\U1/aes_core/SB0/n148 ), .Y(
        \U1/aes_core/SB0/n128 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U47  ( .A0(\U1/aes_core/SB0/n145 ), .A1(
        \U1/aes_core/SB0/n101 ), .B0(\U1/aes_core/SB0/n112 ), .Y(
        \U1/aes_core/SB0/n137 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U46  ( .A0(\U1/aes_core/SB0/n121 ), .A1(
        \U1/aes_core/SB0/n144 ), .B0(\U1/aes_core/SB0/n113 ), .Y(
        \U1/aes_core/SB0/n138 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U45  ( .A0(\U1/aes_core/SB0/n141 ), .A1(
        \U1/aes_core/SB0/n142 ), .B0(\U1/aes_core/SB0/n143 ), .Y(
        \U1/aes_core/SB0/n139 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U44  ( .A(\U1/aes_core/SB0/n137 ), .B(
        \U1/aes_core/SB0/n138 ), .C(\U1/aes_core/SB0/n139 ), .D(
        \U1/aes_core/SB0/n140 ), .Y(\U1/aes_core/SB0/n129 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U43  ( .A(\U1/aes_core/SB0/n106 ), .B(
        \U1/aes_core/SB0/n136 ), .Y(\U1/aes_core/SB0/n104 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB0/U42  ( .A(\U1/aes_core/SB0/n116 ), .B(
        \U1/aes_core/SB0/n104 ), .Y(\U1/aes_core/SB0/n132 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U41  ( .A0(\U1/aes_core/SB0/n118 ), .A1(
        \U1/aes_core/SB0/n131 ), .B0(\U1/aes_core/SB0/n132 ), .B1(
        \U1/aes_core/SB0/n133 ), .C0(\U1/aes_core/SB0/n134 ), .C1(
        \U1/aes_core/SB0/n135 ), .Y(\U1/aes_core/SB0/n130 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U40  ( .A(\U1/aes_core/SB0/n125 ), .B(
        \U1/aes_core/SB0/n126 ), .C(\U1/aes_core/SB0/n127 ), .D(
        \U1/aes_core/SB0/n128 ), .E(\U1/aes_core/SB0/n129 ), .F(
        \U1/aes_core/SB0/n130 ), .Y(\U1/aes_core/sb0 [6]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U39  ( .A0(\U1/aes_core/SB0/n121 ), .A1(
        \U1/aes_core/SB0/n122 ), .B0(\U1/aes_core/SB0/n123 ), .B1(
        \U1/aes_core/SB0/n124 ), .Y(\U1/aes_core/SB0/n120 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB0/U38  ( .A0(\U1/aes_core/SB0/n117 ), .A1(
        \U1/aes_core/SB0/n118 ), .B0(\U1/aes_core/SB0/n119 ), .C0(
        \U1/aes_core/SB0/n120 ), .Y(\U1/aes_core/SB0/n93 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB0/U37  ( .A1N(\U1/aes_core/SB0/n114 ), 
        .A0(\U1/aes_core/SB0/n115 ), .B0(\U1/aes_core/SB0/n116 ), .Y(
        \U1/aes_core/SB0/n107 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U36  ( .A0(\U1/aes_core/SB0/n111 ), .A1(
        \U1/aes_core/SB0/n112 ), .B0(\U1/aes_core/SB0/n113 ), .Y(
        \U1/aes_core/SB0/n108 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U35  ( .A(\U1/aes_core/SB0/n107 ), .B(
        \U1/aes_core/SB0/n108 ), .C(\U1/aes_core/SB0/n109 ), .D(
        \U1/aes_core/SB0/n110 ), .Y(\U1/aes_core/SB0/n94 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U34  ( .A(\U1/aes_core/SB0/n105 ), .B(
        \U1/aes_core/SB0/n106 ), .Y(\U1/aes_core/SB0/n102 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U33  ( .A0(\U1/aes_core/SB0/n101 ), .A1(
        \U1/aes_core/SB0/n102 ), .B0(\U1/aes_core/SB0/n103 ), .B1(
        \U1/aes_core/SB0/n104 ), .Y(\U1/aes_core/SB0/n100 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U32  ( .A0(\U1/aes_core/SB0/n96 ), .A1(
        \U1/aes_core/SB0/n97 ), .B0(\U1/aes_core/SB0/n98 ), .B1(
        \U1/aes_core/SB0/n99 ), .C0(\U1/aes_core/SB0/n100 ), .Y(
        \U1/aes_core/SB0/n95 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U31  ( .A(\U1/aes_core/SB0/n90 ), .B(
        \U1/aes_core/SB0/n91 ), .C(\U1/aes_core/SB0/n92 ), .D(
        \U1/aes_core/SB0/n93 ), .E(\U1/aes_core/SB0/n94 ), .F(
        \U1/aes_core/SB0/n95 ), .Y(\U1/aes_core/sb0 [7]) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U30  ( .A(\U1/aes_core/SB0/n87 ), .B(
        \U1/aes_core/SB0/n88 ), .C(\U1/aes_core/SB0/n89 ), .Y(
        \U1/aes_core/SB0/n64 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U29  ( .A0(\U1/aes_core/SB0/n86 ), .A1(
        \U1/aes_core/SB0/n30 ), .B0(\U1/aes_core/SB0/n14 ), .Y(
        \U1/aes_core/SB0/n81 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U28  ( .A0(\U1/aes_core/SB0/n21 ), .A1(
        \U1/aes_core/SB0/n84 ), .B0(\U1/aes_core/SB0/n85 ), .B1(
        \U1/aes_core/SB0/n20 ), .Y(\U1/aes_core/SB0/n83 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U27  ( .A(\U1/aes_core/SB0/n81 ), .B(
        \U1/aes_core/SB0/n82 ), .C(\U1/aes_core/SB0/n83 ), .Y(
        \U1/aes_core/SB0/n65 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB0/U26  ( .A0(\U1/aes_core/SB0/n78 ), .A1(
        \U1/aes_core/SB0/n55 ), .B0(\U1/aes_core/SB0/n79 ), .B1(
        \U1/aes_core/SB0/n80 ), .Y(\U1/aes_core/SB0/n77 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB0/U25  ( .A0(\U1/aes_core/SB0/n73 ), .A1(
        \U1/aes_core/SB0/n74 ), .B0(\U1/aes_core/SB0/n75 ), .B1(
        \U1/aes_core/SB0/n76 ), .C0(\U1/aes_core/SB0/n77 ), .Y(
        \U1/aes_core/SB0/n66 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U24  ( .A(\U1/aes_core/SB0/n25 ), .B(
        \U1/aes_core/SB0/n72 ), .Y(\U1/aes_core/SB0/n71 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U23  ( .AN(\U1/aes_core/SB0/n68 ), .B(
        \U1/aes_core/SB0/n69 ), .C(\U1/aes_core/SB0/n70 ), .D(
        \U1/aes_core/SB0/n71 ), .Y(\U1/aes_core/SB0/n67 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U22  ( .A(\U1/aes_core/SB0/n62 ), .B(
        \U1/aes_core/SB0/n63 ), .C(\U1/aes_core/SB0/n64 ), .D(
        \U1/aes_core/SB0/n65 ), .E(\U1/aes_core/SB0/n66 ), .F(
        \U1/aes_core/SB0/n67 ), .Y(\U1/aes_core/SB0/n3 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB0/U21  ( .A(\U1/aes_core/SB0/n59 ), .B(
        \U1/aes_core/SB0/n60 ), .C(\U1/aes_core/SB0/n61 ), .D(
        \U1/aes_core/SB0/n3 ), .Y(\U1/aes_core/SB0/n34 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U20  ( .A0(\U1/aes_core/SB0/n57 ), .A1(
        \U1/aes_core/SB0/n46 ), .B0(\U1/aes_core/SB0/n10 ), .B1(
        \U1/aes_core/SB0/n58 ), .Y(\U1/aes_core/SB0/n56 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U19  ( .A0(\U1/aes_core/SB0/n32 ), .A1(
        \U1/aes_core/SB0/n20 ), .B0(\U1/aes_core/SB0/n29 ), .B1(
        \U1/aes_core/SB0/n55 ), .C0(\U1/aes_core/SB0/n56 ), .Y(
        \U1/aes_core/SB0/n35 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB0/U18  ( .A0(\U1/aes_core/SB0/n51 ), .A1(
        \U1/aes_core/SB0/n52 ), .B0(\U1/aes_core/SB0/n53 ), .B1(
        \U1/aes_core/SB0/n54 ), .Y(\U1/aes_core/SB0/n50 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U17  ( .A0(\U1/aes_core/SB0/n47 ), .A1(
        \U1/aes_core/SB0/n48 ), .B0(\U1/aes_core/SB0/n49 ), .B1(
        \U1/aes_core/SB0/n24 ), .C0(\U1/aes_core/SB0/n50 ), .Y(
        \U1/aes_core/SB0/n36 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB0/U16  ( .A(\U1/aes_core/SB0/n45 ), .B(
        \U1/aes_core/SB0/n46 ), .Y(\U1/aes_core/SB0/n38 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U15  ( .A(\U1/aes_core/SB0/n44 ), .Y(
        \U1/aes_core/SB0/n39 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB0/U14  ( .A(\U1/aes_core/SB0/n41 ), .B(
        \U1/aes_core/SB0/n42 ), .C(\U1/aes_core/SB0/n43 ), .Y(
        \U1/aes_core/SB0/n40 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U13  ( .A0(\U1/aes_core/SB0/n23 ), .A1(
        \U1/aes_core/SB0/n38 ), .B0(\U1/aes_core/SB0/n31 ), .B1(
        \U1/aes_core/SB0/n39 ), .C0(\U1/aes_core/SB0/n40 ), .Y(
        \U1/aes_core/SB0/n37 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB0/U12  ( .AN(\U1/aes_core/SB0/n34 ), .B(
        \U1/aes_core/SB0/n35 ), .C(\U1/aes_core/SB0/n36 ), .D(
        \U1/aes_core/SB0/n37 ), .Y(\U1/aes_core/sb0 [8]) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB0/U11  ( .A0(\U1/aes_core/SB0/n29 ), .A1(
        \U1/aes_core/SB0/n30 ), .B0(\U1/aes_core/SB0/n31 ), .B1(
        \U1/aes_core/SB0/n32 ), .C0(\U1/aes_core/SB0/n33 ), .Y(
        \U1/aes_core/SB0/n28 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB0/U10  ( .A(\U1/aes_core/SB0/n28 ), .Y(
        \U1/aes_core/SB0/n4 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U9  ( .A0(\U1/aes_core/SB0/n15 ), .A1(
        \U1/aes_core/SB0/n26 ), .B0(\U1/aes_core/SB0/n27 ), .Y(
        \U1/aes_core/SB0/n16 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U8  ( .A0(\U1/aes_core/SB0/n23 ), .A1(
        \U1/aes_core/SB0/n24 ), .B0(\U1/aes_core/SB0/n25 ), .Y(
        \U1/aes_core/SB0/n17 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB0/U7  ( .A0(\U1/aes_core/SB0/n20 ), .A1(
        \U1/aes_core/SB0/n21 ), .B0(\U1/aes_core/SB0/n22 ), .Y(
        \U1/aes_core/SB0/n18 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB0/U6  ( .A(\U1/aes_core/SB0/n16 ), .B(
        \U1/aes_core/SB0/n17 ), .C(\U1/aes_core/SB0/n18 ), .D(
        \U1/aes_core/SB0/n19 ), .Y(\U1/aes_core/SB0/n5 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB0/U5  ( .A(\U1/aes_core/SB0/n13 ), .B(
        \U1/aes_core/SB0/n14 ), .C(\U1/aes_core/SB0/n15 ), .Y(
        \U1/aes_core/SB0/n9 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB0/U4  ( .A0(\U1/aes_core/SB0/n7 ), .A1(
        \U1/aes_core/SB0/n8 ), .B0(\U1/aes_core/SB0/n9 ), .B1(
        \U1/aes_core/SB0/n10 ), .C0(\U1/aes_core/SB0/n11 ), .C1(
        \U1/aes_core/SB0/n12 ), .Y(\U1/aes_core/SB0/n6 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB0/U3  ( .A(\U1/aes_core/SB0/n1 ), .B(
        \U1/aes_core/SB0/n2 ), .C(\U1/aes_core/SB0/n3 ), .D(
        \U1/aes_core/SB0/n4 ), .E(\U1/aes_core/SB0/n5 ), .F(
        \U1/aes_core/SB0/n6 ), .Y(\U1/aes_core/sb0 [9]) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U711  ( .A0(\U1/aes_core/SB1/n2402 ), .A1(
        \U1/aes_core/SB1/n2157 ), .B0(\U1/aes_core/SB1/n2480 ), .B1(
        \U1/aes_core/SB1/n2464 ), .C0(\U1/aes_core/SB1/n2225 ), .Y(
        \U1/aes_core/SB1/n2158 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U393  ( .A0(\U1/aes_core/SB1/n2650 ), .A1(
        \U1/aes_core/SB1/n2775 ), .B0(\U1/aes_core/SB1/n2773 ), .B1(
        \U1/aes_core/SB1/n2758 ), .C0(\U1/aes_core/SB1/n2649 ), .Y(
        \U1/aes_core/SB1/n2652 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U391  ( .A0(\U1/aes_core/SB1/n2971 ), .A1(
        \U1/aes_core/SB1/n3096 ), .B0(\U1/aes_core/SB1/n3094 ), .B1(
        \U1/aes_core/SB1/n3079 ), .C0(\U1/aes_core/SB1/n2970 ), .Y(
        \U1/aes_core/SB1/n2973 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U363  ( .A0(\U1/aes_core/SB1/n2203 ), .A1(
        \U1/aes_core/SB1/n2353 ), .B0(\U1/aes_core/SB1/n2351 ), .B1(
        \U1/aes_core/SB1/n2311 ), .C0(\U1/aes_core/SB1/n2202 ), .Y(
        \U1/aes_core/SB1/n2205 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U361  ( .A0(\U1/aes_core/SB1/n2824 ), .A1(
        \U1/aes_core/SB1/n2604 ), .B0(\U1/aes_core/SB1/n2923 ), .B1(
        \U1/aes_core/SB1/n2907 ), .C0(\U1/aes_core/SB1/n2672 ), .Y(
        \U1/aes_core/SB1/n2605 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U301  ( .A0(\U1/aes_core/SB1/n3145 ), .A1(
        \U1/aes_core/SB1/n2328 ), .B0(\U1/aes_core/SB1/n3223 ), .B1(
        \U1/aes_core/SB1/n3207 ), .C0(\U1/aes_core/SB1/n2993 ), .Y(
        \U1/aes_core/SB1/n2329 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U300  ( .A0(\U1/aes_core/SB1/n2402 ), .A1(
        \U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2480 ), .B1(
        \U1/aes_core/SB1/n2478 ), .C0(\U1/aes_core/SB1/n2268 ), .Y(
        \U1/aes_core/SB1/n2144 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U151  ( .A0(\U1/aes_core/SB1/n2824 ), .A1(
        \U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2923 ), .B1(
        \U1/aes_core/SB1/n2921 ), .C0(\U1/aes_core/SB1/n2715 ), .Y(
        \U1/aes_core/SB1/n2591 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB1/U150  ( .A0(\U1/aes_core/SB1/n3145 ), .A1(
        \U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3223 ), .B1(
        \U1/aes_core/SB1/n3221 ), .C0(\U1/aes_core/SB1/n3036 ), .Y(
        \U1/aes_core/SB1/n1742 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1724  ( .A(Dout[71]), .B(Dout[70]), .Y(
        \U1/aes_core/SB1/n1691 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1723  ( .A(Dout[69]), .B(Dout[68]), .Y(
        \U1/aes_core/SB1/n1682 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1722  ( .A(\U1/aes_core/SB1/n1691 ), .B(
        \U1/aes_core/SB1/n1682 ), .Y(\U1/aes_core/SB1/n2328 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1721  ( .A(Dout[65]), .Y(
        \U1/aes_core/SB1/n767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1720  ( .A(Dout[64]), .Y(
        \U1/aes_core/SB1/n385 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1719  ( .A(\U1/aes_core/SB1/n767 ), .B(
        \U1/aes_core/SB1/n385 ), .Y(\U1/aes_core/SB1/n1683 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1718  ( .A(Dout[67]), .B(Dout[66]), .Y(
        \U1/aes_core/SB1/n1703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1717  ( .A(\U1/aes_core/SB1/n1683 ), .B(
        \U1/aes_core/SB1/n1703 ), .Y(\U1/aes_core/SB1/n3207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1716  ( .A(\U1/aes_core/SB1/n2328 ), .B(
        \U1/aes_core/SB1/n3207 ), .Y(\U1/aes_core/SB1/n3014 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U1715  ( .A(Dout[66]), .B(Dout[67]), .Y(
        \U1/aes_core/SB1/n1686 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1714  ( .A(\U1/aes_core/SB1/n1686 ), .B(
        \U1/aes_core/SB1/n1683 ), .Y(\U1/aes_core/SB1/n3145 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1713  ( .A(Dout[71]), .Y(
        \U1/aes_core/SB1/n1203 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1712  ( .A(\U1/aes_core/SB1/n1203 ), .B(
        Dout[70]), .Y(\U1/aes_core/SB1/n1709 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1711  ( .A(\U1/aes_core/SB1/n1709 ), .B(
        \U1/aes_core/SB1/n1682 ), .Y(\U1/aes_core/SB1/n2327 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1710  ( .A(\U1/aes_core/SB1/n3145 ), .B(
        \U1/aes_core/SB1/n2327 ), .Y(\U1/aes_core/SB1/n3111 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1709  ( .A(Dout[67]), .Y(
        \U1/aes_core/SB1/n707 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U1708  ( .A(Dout[66]), .B(
        \U1/aes_core/SB1/n707 ), .Y(\U1/aes_core/SB1/n1684 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1707  ( .A(\U1/aes_core/SB1/n1683 ), .B(
        \U1/aes_core/SB1/n1684 ), .Y(\U1/aes_core/SB1/n3076 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1706  ( .A(\U1/aes_core/SB1/n3076 ), .Y(
        \U1/aes_core/SB1/n3241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1705  ( .A(Dout[68]), .Y(
        \U1/aes_core/SB1/n752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1704  ( .A(\U1/aes_core/SB1/n752 ), .B(
        Dout[69]), .Y(\U1/aes_core/SB1/n1690 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1703  ( .A(Dout[70]), .Y(
        \U1/aes_core/SB1/n1158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1702  ( .A(\U1/aes_core/SB1/n1158 ), .B(
        Dout[71]), .Y(\U1/aes_core/SB1/n1700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1701  ( .A(\U1/aes_core/SB1/n1690 ), .B(
        \U1/aes_core/SB1/n1700 ), .Y(\U1/aes_core/SB1/n3097 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1700  ( .A(\U1/aes_core/SB1/n3097 ), .Y(
        \U1/aes_core/SB1/n3195 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1699  ( .A(\U1/aes_core/SB1/n3241 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n3054 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1698  ( .A(\U1/aes_core/SB1/n2328 ), .Y(
        \U1/aes_core/SB1/n3210 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1697  ( .A(Dout[65]), .B(Dout[64]), .Y(
        \U1/aes_core/SB1/n1687 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1696  ( .A(\U1/aes_core/SB1/n1687 ), .B(
        \U1/aes_core/SB1/n1703 ), .Y(\U1/aes_core/SB1/n3163 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1695  ( .A(\U1/aes_core/SB1/n3163 ), .Y(
        \U1/aes_core/SB1/n3251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1694  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3251 ), .Y(\U1/aes_core/SB1/n3168 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1693  ( .A(\U1/aes_core/SB1/n385 ), .B(
        Dout[65]), .Y(\U1/aes_core/SB1/n1702 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1692  ( .A(\U1/aes_core/SB1/n1684 ), .B(
        \U1/aes_core/SB1/n1702 ), .Y(\U1/aes_core/SB1/n3063 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1691  ( .A(\U1/aes_core/SB1/n3063 ), .Y(
        \U1/aes_core/SB1/n3152 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1690  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3032 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U1689  ( .A(\U1/aes_core/SB1/n3054 ), .B(
        \U1/aes_core/SB1/n3168 ), .C(\U1/aes_core/SB1/n3032 ), .Y(
        \U1/aes_core/SB1/n1722 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1688  ( .A(\U1/aes_core/SB1/n1682 ), .B(
        \U1/aes_core/SB1/n1700 ), .Y(\U1/aes_core/SB1/n3096 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1687  ( .A(\U1/aes_core/SB1/n707 ), .B(
        Dout[66]), .Y(\U1/aes_core/SB1/n1693 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1686  ( .A(\U1/aes_core/SB1/n1693 ), .B(
        \U1/aes_core/SB1/n1702 ), .Y(\U1/aes_core/SB1/n3094 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1685  ( .A(\U1/aes_core/SB1/n3096 ), .B(
        \U1/aes_core/SB1/n3094 ), .Y(\U1/aes_core/SB1/n3009 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1684  ( .A(\U1/aes_core/SB1/n2327 ), .Y(
        \U1/aes_core/SB1/n3212 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1683  ( .A(Dout[69]), .Y(
        \U1/aes_core/SB1/n1030 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1682  ( .A(\U1/aes_core/SB1/n752 ), .B(
        \U1/aes_core/SB1/n1030 ), .Y(\U1/aes_core/SB1/n1701 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1681  ( .A(\U1/aes_core/SB1/n1691 ), .B(
        \U1/aes_core/SB1/n1701 ), .Y(\U1/aes_core/SB1/n3255 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1680  ( .A(\U1/aes_core/SB1/n3255 ), .Y(
        \U1/aes_core/SB1/n3186 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1679  ( .A(\U1/aes_core/SB1/n767 ), .B(
        Dout[64]), .Y(\U1/aes_core/SB1/n1692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1678  ( .A(\U1/aes_core/SB1/n1692 ), .B(
        \U1/aes_core/SB1/n1703 ), .Y(\U1/aes_core/SB1/n3220 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1677  ( .A(\U1/aes_core/SB1/n3220 ), .Y(
        \U1/aes_core/SB1/n3068 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1676  ( .A0(\U1/aes_core/SB1/n3212 ), 
        .A1(\U1/aes_core/SB1/n3186 ), .B0(\U1/aes_core/SB1/n3068 ), .Y(
        \U1/aes_core/SB1/n1621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1675  ( .A(\U1/aes_core/SB1/n1687 ), .B(
        \U1/aes_core/SB1/n1684 ), .Y(\U1/aes_core/SB1/n3208 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1674  ( .A(\U1/aes_core/SB1/n3208 ), .Y(
        \U1/aes_core/SB1/n3194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1673  ( .A(\U1/aes_core/SB1/n1030 ), .B(
        Dout[68]), .Y(\U1/aes_core/SB1/n1708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1672  ( .A(\U1/aes_core/SB1/n1700 ), .B(
        \U1/aes_core/SB1/n1708 ), .Y(\U1/aes_core/SB1/n3248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1671  ( .A(\U1/aes_core/SB1/n3096 ), .B(
        \U1/aes_core/SB1/n3248 ), .Y(\U1/aes_core/SB1/n2987 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1670  ( .A(\U1/aes_core/SB1/n1203 ), .B(
        \U1/aes_core/SB1/n1158 ), .Y(\U1/aes_core/SB1/n1699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1669  ( .A(\U1/aes_core/SB1/n1690 ), .B(
        \U1/aes_core/SB1/n1699 ), .Y(\U1/aes_core/SB1/n3223 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1668  ( .A(\U1/aes_core/SB1/n3223 ), .Y(
        \U1/aes_core/SB1/n2968 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1667  ( .A0(\U1/aes_core/SB1/n3194 ), 
        .A1(\U1/aes_core/SB1/n2987 ), .B0(\U1/aes_core/SB1/n2968 ), .B1(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n1218 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1666  ( .AN(\U1/aes_core/SB1/n3009 ), 
        .B(\U1/aes_core/SB1/n1621 ), .C(\U1/aes_core/SB1/n1218 ), .Y(
        \U1/aes_core/SB1/n1721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1665  ( .A(\U1/aes_core/SB1/n1682 ), .B(
        \U1/aes_core/SB1/n1699 ), .Y(\U1/aes_core/SB1/n3113 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1664  ( .A(\U1/aes_core/SB1/n1686 ), .B(
        \U1/aes_core/SB1/n1687 ), .Y(\U1/aes_core/SB1/n3258 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1663  ( .A(\U1/aes_core/SB1/n1709 ), .B(
        \U1/aes_core/SB1/n1690 ), .Y(\U1/aes_core/SB1/n3164 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1662  ( .A(\U1/aes_core/SB1/n1686 ), .B(
        \U1/aes_core/SB1/n1692 ), .Y(\U1/aes_core/SB1/n3161 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1661  ( .A(\U1/aes_core/SB1/n1683 ), .B(
        \U1/aes_core/SB1/n1693 ), .Y(\U1/aes_core/SB1/n3166 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1660  ( .A(\U1/aes_core/SB1/n3166 ), .Y(
        \U1/aes_core/SB1/n3146 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1659  ( .A(\U1/aes_core/SB1/n3248 ), .Y(
        \U1/aes_core/SB1/n2982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1658  ( .A(\U1/aes_core/SB1/n1684 ), .B(
        \U1/aes_core/SB1/n1692 ), .Y(\U1/aes_core/SB1/n3184 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1657  ( .A(\U1/aes_core/SB1/n3184 ), .Y(
        \U1/aes_core/SB1/n3209 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1656  ( .A0(\U1/aes_core/SB1/n3146 ), 
        .A1(\U1/aes_core/SB1/n3210 ), .B0(\U1/aes_core/SB1/n2982 ), .B1(
        \U1/aes_core/SB1/n3209 ), .Y(\U1/aes_core/SB1/n1685 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1655  ( .A0(\U1/aes_core/SB1/n3113 ), 
        .A1(\U1/aes_core/SB1/n3258 ), .B0(\U1/aes_core/SB1/n3164 ), .B1(
        \U1/aes_core/SB1/n3161 ), .C0(\U1/aes_core/SB1/n1685 ), .Y(
        \U1/aes_core/SB1/n1720 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1654  ( .A(\U1/aes_core/SB1/n3166 ), .B(
        \U1/aes_core/SB1/n3113 ), .Y(\U1/aes_core/SB1/n2975 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1653  ( .A(\U1/aes_core/SB1/n3161 ), .B(
        \U1/aes_core/SB1/n3096 ), .Y(\U1/aes_core/SB1/n2985 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1652  ( .A(\U1/aes_core/SB1/n2985 ), .Y(
        \U1/aes_core/SB1/n1689 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1651  ( .A(\U1/aes_core/SB1/n1686 ), .B(
        \U1/aes_core/SB1/n1702 ), .Y(\U1/aes_core/SB1/n3236 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1650  ( .A(\U1/aes_core/SB1/n3236 ), .Y(
        \U1/aes_core/SB1/n3185 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1649  ( .A(\U1/aes_core/SB1/n1687 ), .B(
        \U1/aes_core/SB1/n1693 ), .Y(\U1/aes_core/SB1/n3221 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1648  ( .A(\U1/aes_core/SB1/n3221 ), .Y(
        \U1/aes_core/SB1/n3232 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1647  ( .A0(\U1/aes_core/SB1/n3185 ), 
        .A1(\U1/aes_core/SB1/n3232 ), .B0(\U1/aes_core/SB1/n3186 ), .Y(
        \U1/aes_core/SB1/n1688 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1646  ( .A(\U1/aes_core/SB1/n1691 ), .B(
        \U1/aes_core/SB1/n1708 ), .Y(\U1/aes_core/SB1/n3237 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1645  ( .A(\U1/aes_core/SB1/n3237 ), .Y(
        \U1/aes_core/SB1/n3187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1644  ( .A(\U1/aes_core/SB1/n3187 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3002 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1643  ( .AN(\U1/aes_core/SB1/n2975 ), 
        .B(\U1/aes_core/SB1/n1689 ), .C(\U1/aes_core/SB1/n1688 ), .D(
        \U1/aes_core/SB1/n3002 ), .Y(\U1/aes_core/SB1/n1698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1642  ( .A(\U1/aes_core/SB1/n1701 ), .B(
        \U1/aes_core/SB1/n1699 ), .Y(\U1/aes_core/SB1/n3257 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1641  ( .A(\U1/aes_core/SB1/n1691 ), .B(
        \U1/aes_core/SB1/n1690 ), .Y(\U1/aes_core/SB1/n3249 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1640  ( .A0(\U1/aes_core/SB1/n2327 ), 
        .A1(\U1/aes_core/SB1/n3076 ), .B0(\U1/aes_core/SB1/n3257 ), .B1(
        \U1/aes_core/SB1/n3166 ), .C0(\U1/aes_core/SB1/n3249 ), .C1(
        \U1/aes_core/SB1/n3184 ), .Y(\U1/aes_core/SB1/n1697 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1639  ( .A(\U1/aes_core/SB1/n3208 ), .B(
        \U1/aes_core/SB1/n2327 ), .Y(\U1/aes_core/SB1/n3060 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1638  ( .A(\U1/aes_core/SB1/n2982 ), .B(
        \U1/aes_core/SB1/n3146 ), .Y(\U1/aes_core/SB1/n3013 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1637  ( .A(\U1/aes_core/SB1/n3209 ), .B(
        \U1/aes_core/SB1/n3210 ), .Y(\U1/aes_core/SB1/n3033 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1636  ( .A(\U1/aes_core/SB1/n3164 ), .Y(
        \U1/aes_core/SB1/n3238 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1635  ( .A(\U1/aes_core/SB1/n3238 ), .B(
        \U1/aes_core/SB1/n3068 ), .Y(\U1/aes_core/SB1/n3071 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1634  ( .AN(\U1/aes_core/SB1/n3060 ), 
        .B(\U1/aes_core/SB1/n3013 ), .C(\U1/aes_core/SB1/n3033 ), .D(
        \U1/aes_core/SB1/n3071 ), .Y(\U1/aes_core/SB1/n1696 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1633  ( .A(\U1/aes_core/SB1/n1709 ), .B(
        \U1/aes_core/SB1/n1701 ), .Y(\U1/aes_core/SB1/n2983 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1632  ( .A(\U1/aes_core/SB1/n2983 ), .B(
        \U1/aes_core/SB1/n3220 ), .Y(\U1/aes_core/SB1/n3137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1631  ( .A(\U1/aes_core/SB1/n1693 ), .B(
        \U1/aes_core/SB1/n1692 ), .Y(\U1/aes_core/SB1/n3256 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1630  ( .A(\U1/aes_core/SB1/n3223 ), .B(
        \U1/aes_core/SB1/n3256 ), .Y(\U1/aes_core/SB1/n3102 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1629  ( .A(\U1/aes_core/SB1/n3102 ), .Y(
        \U1/aes_core/SB1/n1694 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1628  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3068 ), .Y(\U1/aes_core/SB1/n3121 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1627  ( .A(\U1/aes_core/SB1/n3256 ), .Y(
        \U1/aes_core/SB1/n3239 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1626  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3239 ), .Y(\U1/aes_core/SB1/n3172 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1625  ( .AN(\U1/aes_core/SB1/n3137 ), 
        .B(\U1/aes_core/SB1/n1694 ), .C(\U1/aes_core/SB1/n3121 ), .D(
        \U1/aes_core/SB1/n3172 ), .Y(\U1/aes_core/SB1/n1695 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1624  ( .A(\U1/aes_core/SB1/n1698 ), .B(
        \U1/aes_core/SB1/n1697 ), .C(\U1/aes_core/SB1/n1696 ), .D(
        \U1/aes_core/SB1/n1695 ), .Y(\U1/aes_core/SB1/n2905 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1623  ( .A(\U1/aes_core/SB1/n3163 ), .B(
        \U1/aes_core/SB1/n2983 ), .Y(\U1/aes_core/SB1/n3171 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1622  ( .A(\U1/aes_core/SB1/n1708 ), .B(
        \U1/aes_core/SB1/n1699 ), .Y(\U1/aes_core/SB1/n3079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1621  ( .A(\U1/aes_core/SB1/n3145 ), .B(
        \U1/aes_core/SB1/n3079 ), .Y(\U1/aes_core/SB1/n3050 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1620  ( .A(\U1/aes_core/SB1/n3257 ), .Y(
        \U1/aes_core/SB1/n3213 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1619  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3194 ), .Y(\U1/aes_core/SB1/n2999 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1618  ( .A0(\U1/aes_core/SB1/n3079 ), 
        .A1(\U1/aes_core/SB1/n3256 ), .B0(\U1/aes_core/SB1/n2999 ), .Y(
        \U1/aes_core/SB1/n1707 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1617  ( .A(\U1/aes_core/SB1/n3094 ), .Y(
        \U1/aes_core/SB1/n3189 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1616  ( .A(\U1/aes_core/SB1/n3189 ), .B(
        \U1/aes_core/SB1/n3212 ), .Y(\U1/aes_core/SB1/n3190 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1615  ( .A(\U1/aes_core/SB1/n3212 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1614  ( .A(\U1/aes_core/SB1/n1701 ), .B(
        \U1/aes_core/SB1/n1700 ), .Y(\U1/aes_core/SB1/n3219 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1613  ( .A(\U1/aes_core/SB1/n3219 ), .Y(
        \U1/aes_core/SB1/n2994 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1612  ( .A(\U1/aes_core/SB1/n3185 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3018 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1611  ( .A(\U1/aes_core/SB1/n3207 ), .Y(
        \U1/aes_core/SB1/n3188 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1610  ( .A(\U1/aes_core/SB1/n3188 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3082 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1609  ( .A(\U1/aes_core/SB1/n3190 ), .B(
        \U1/aes_core/SB1/n3149 ), .C(\U1/aes_core/SB1/n3018 ), .D(
        \U1/aes_core/SB1/n3082 ), .Y(\U1/aes_core/SB1/n1706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1608  ( .A(\U1/aes_core/SB1/n3209 ), .B(
        \U1/aes_core/SB1/n3187 ), .Y(\U1/aes_core/SB1/n3116 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1607  ( .A(\U1/aes_core/SB1/n3251 ), .B(
        \U1/aes_core/SB1/n3187 ), .Y(\U1/aes_core/SB1/n3107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1606  ( .A(\U1/aes_core/SB1/n3249 ), .Y(
        \U1/aes_core/SB1/n3242 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1605  ( .A(\U1/aes_core/SB1/n3146 ), .B(
        \U1/aes_core/SB1/n3242 ), .Y(\U1/aes_core/SB1/n2979 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1604  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3185 ), .Y(\U1/aes_core/SB1/n3090 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1603  ( .A(\U1/aes_core/SB1/n3116 ), .B(
        \U1/aes_core/SB1/n3107 ), .C(\U1/aes_core/SB1/n2979 ), .D(
        \U1/aes_core/SB1/n3090 ), .Y(\U1/aes_core/SB1/n1705 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1602  ( .A(\U1/aes_core/SB1/n3161 ), .Y(
        \U1/aes_core/SB1/n3130 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1601  ( .A(\U1/aes_core/SB1/n2982 ), .B(
        \U1/aes_core/SB1/n3130 ), .Y(\U1/aes_core/SB1/n2966 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1600  ( .A(\U1/aes_core/SB1/n1703 ), .B(
        \U1/aes_core/SB1/n1702 ), .Y(\U1/aes_core/SB1/n3196 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1599  ( .A(\U1/aes_core/SB1/n3196 ), .Y(
        \U1/aes_core/SB1/n3230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1598  ( .A(\U1/aes_core/SB1/n2982 ), .B(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n3030 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1597  ( .A(\U1/aes_core/SB1/n3145 ), .Y(
        \U1/aes_core/SB1/n3253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1596  ( .A(\U1/aes_core/SB1/n3253 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n3065 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1595  ( .A(\U1/aes_core/SB1/n3186 ), .B(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n3214 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1594  ( .A(\U1/aes_core/SB1/n2966 ), .B(
        \U1/aes_core/SB1/n3030 ), .C(\U1/aes_core/SB1/n3065 ), .D(
        \U1/aes_core/SB1/n3214 ), .Y(\U1/aes_core/SB1/n1704 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1593  ( .A(\U1/aes_core/SB1/n3171 ), .B(
        \U1/aes_core/SB1/n3050 ), .C(\U1/aes_core/SB1/n1707 ), .D(
        \U1/aes_core/SB1/n1706 ), .E(\U1/aes_core/SB1/n1705 ), .F(
        \U1/aes_core/SB1/n1704 ), .Y(\U1/aes_core/SB1/n2894 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1592  ( .A(\U1/aes_core/SB1/n2894 ), .Y(
        \U1/aes_core/SB1/n1718 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1591  ( .A(\U1/aes_core/SB1/n3221 ), .B(
        \U1/aes_core/SB1/n3079 ), .Y(\U1/aes_core/SB1/n2976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1590  ( .A(\U1/aes_core/SB1/n1709 ), .B(
        \U1/aes_core/SB1/n1708 ), .Y(\U1/aes_core/SB1/n3218 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1589  ( .A(\U1/aes_core/SB1/n3218 ), .B(
        \U1/aes_core/SB1/n3094 ), .Y(\U1/aes_core/SB1/n3103 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1588  ( .A(\U1/aes_core/SB1/n3103 ), .Y(
        \U1/aes_core/SB1/n1711 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1587  ( .A(\U1/aes_core/SB1/n3096 ), .Y(
        \U1/aes_core/SB1/n3243 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1586  ( .A0(\U1/aes_core/SB1/n2994 ), 
        .A1(\U1/aes_core/SB1/n3243 ), .B0(\U1/aes_core/SB1/n3230 ), .Y(
        \U1/aes_core/SB1/n1710 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1585  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3130 ), .Y(\U1/aes_core/SB1/n3001 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1584  ( .AN(\U1/aes_core/SB1/n2976 ), 
        .B(\U1/aes_core/SB1/n1711 ), .C(\U1/aes_core/SB1/n1710 ), .D(
        \U1/aes_core/SB1/n3001 ), .Y(\U1/aes_core/SB1/n1715 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1583  ( .A0(\U1/aes_core/SB1/n3207 ), 
        .A1(\U1/aes_core/SB1/n3255 ), .B0(\U1/aes_core/SB1/n3113 ), .B1(
        \U1/aes_core/SB1/n3161 ), .C0(\U1/aes_core/SB1/n3220 ), .C1(
        \U1/aes_core/SB1/n3237 ), .Y(\U1/aes_core/SB1/n1714 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1582  ( .A(\U1/aes_core/SB1/n3255 ), .B(
        \U1/aes_core/SB1/n3258 ), .Y(\U1/aes_core/SB1/n3041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1581  ( .A(\U1/aes_core/SB1/n3243 ), .B(
        \U1/aes_core/SB1/n3185 ), .Y(\U1/aes_core/SB1/n3174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1580  ( .A(\U1/aes_core/SB1/n3146 ), .B(
        \U1/aes_core/SB1/n3243 ), .Y(\U1/aes_core/SB1/n3108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1579  ( .A(\U1/aes_core/SB1/n3130 ), .B(
        \U1/aes_core/SB1/n3210 ), .Y(\U1/aes_core/SB1/n2980 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1578  ( .AN(\U1/aes_core/SB1/n3041 ), 
        .B(\U1/aes_core/SB1/n3174 ), .C(\U1/aes_core/SB1/n3108 ), .D(
        \U1/aes_core/SB1/n2980 ), .Y(\U1/aes_core/SB1/n1713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1577  ( .A(\U1/aes_core/SB1/n3253 ), .B(
        \U1/aes_core/SB1/n3238 ), .Y(\U1/aes_core/SB1/n3053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1576  ( .A(\U1/aes_core/SB1/n3130 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3120 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1575  ( .A(\U1/aes_core/SB1/n2982 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3021 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1574  ( .A(\U1/aes_core/SB1/n3189 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n3066 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1573  ( .A(\U1/aes_core/SB1/n3053 ), .B(
        \U1/aes_core/SB1/n3120 ), .C(\U1/aes_core/SB1/n3021 ), .D(
        \U1/aes_core/SB1/n3066 ), .Y(\U1/aes_core/SB1/n1712 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1572  ( .A(\U1/aes_core/SB1/n1715 ), .B(
        \U1/aes_core/SB1/n1714 ), .C(\U1/aes_core/SB1/n1713 ), .D(
        \U1/aes_core/SB1/n1712 ), .Y(\U1/aes_core/SB1/n1716 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1571  ( .A(\U1/aes_core/SB1/n1716 ), .Y(
        \U1/aes_core/SB1/n3235 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1570  ( .A(\U1/aes_core/SB1/n3251 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n1717 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1569  ( .AN(\U1/aes_core/SB1/n2905 ), 
        .B(\U1/aes_core/SB1/n1718 ), .C(\U1/aes_core/SB1/n3235 ), .D(
        \U1/aes_core/SB1/n1717 ), .Y(\U1/aes_core/SB1/n1719 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1568  ( .A(\U1/aes_core/SB1/n3014 ), .B(
        \U1/aes_core/SB1/n3111 ), .C(\U1/aes_core/SB1/n1722 ), .D(
        \U1/aes_core/SB1/n1721 ), .E(\U1/aes_core/SB1/n1720 ), .F(
        \U1/aes_core/SB1/n1719 ), .Y(\U1/aes_core/SB1/n2346 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1567  ( .A(\U1/aes_core/SB1/n3236 ), .B(
        \U1/aes_core/SB1/n2327 ), .Y(\U1/aes_core/SB1/n3059 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1566  ( .A(\U1/aes_core/SB1/n3186 ), .B(
        \U1/aes_core/SB1/n3253 ), .Y(\U1/aes_core/SB1/n3110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1565  ( .A(\U1/aes_core/SB1/n3242 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3012 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1564  ( .A(\U1/aes_core/SB1/n2983 ), .Y(
        \U1/aes_core/SB1/n3231 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1563  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3035 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1562  ( .AN(\U1/aes_core/SB1/n3059 ), 
        .B(\U1/aes_core/SB1/n3110 ), .C(\U1/aes_core/SB1/n3012 ), .D(
        \U1/aes_core/SB1/n3035 ), .Y(\U1/aes_core/SB1/n1729 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1561  ( .A(\U1/aes_core/SB1/n3223 ), .B(
        \U1/aes_core/SB1/n3094 ), .Y(\U1/aes_core/SB1/n3136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1560  ( .A(\U1/aes_core/SB1/n3146 ), .B(
        \U1/aes_core/SB1/n3212 ), .Y(\U1/aes_core/SB1/n2992 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1559  ( .A0(\U1/aes_core/SB1/n3232 ), 
        .A1(\U1/aes_core/SB1/n3152 ), .B0(\U1/aes_core/SB1/n2982 ), .Y(
        \U1/aes_core/SB1/n1723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1558  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3084 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1557  ( .AN(\U1/aes_core/SB1/n3136 ), 
        .B(\U1/aes_core/SB1/n2992 ), .C(\U1/aes_core/SB1/n1723 ), .D(
        \U1/aes_core/SB1/n3084 ), .Y(\U1/aes_core/SB1/n1724 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1556  ( .A(\U1/aes_core/SB1/n1724 ), .Y(
        \U1/aes_core/SB1/n1728 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1555  ( .A(\U1/aes_core/SB1/n3113 ), .Y(
        \U1/aes_core/SB1/n3233 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1554  ( .A(\U1/aes_core/SB1/n3258 ), .Y(
        \U1/aes_core/SB1/n3153 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U1553  ( .A0(\U1/aes_core/SB1/n3253 ), 
        .A1(\U1/aes_core/SB1/n3187 ), .B0(\U1/aes_core/SB1/n3233 ), .B1(
        \U1/aes_core/SB1/n3068 ), .C0(\U1/aes_core/SB1/n3153 ), .C1(
        \U1/aes_core/SB1/n3231 ), .Y(\U1/aes_core/SB1/n1727 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1552  ( .A0(\U1/aes_core/SB1/n3079 ), 
        .A1(\U1/aes_core/SB1/n3236 ), .B0(\U1/aes_core/SB1/n3256 ), .B1(
        \U1/aes_core/SB1/n3257 ), .Y(\U1/aes_core/SB1/n1725 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1551  ( .A0(\U1/aes_core/SB1/n3130 ), 
        .A1(\U1/aes_core/SB1/n2968 ), .B0(\U1/aes_core/SB1/n3186 ), .B1(
        \U1/aes_core/SB1/n3209 ), .C0(\U1/aes_core/SB1/n1725 ), .Y(
        \U1/aes_core/SB1/n1726 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1550  ( .AN(\U1/aes_core/SB1/n1729 ), 
        .B(\U1/aes_core/SB1/n1728 ), .C(\U1/aes_core/SB1/n1727 ), .D(
        \U1/aes_core/SB1/n1726 ), .Y(\U1/aes_core/SB1/n2903 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1549  ( .A(\U1/aes_core/SB1/n3257 ), .B(
        \U1/aes_core/SB1/n3094 ), .Y(\U1/aes_core/SB1/n2977 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1548  ( .A0(\U1/aes_core/SB1/n3164 ), 
        .A1(\U1/aes_core/SB1/n3257 ), .B0(\U1/aes_core/SB1/n3196 ), .Y(
        \U1/aes_core/SB1/n1734 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1547  ( .A(\U1/aes_core/SB1/n3196 ), .B(
        \U1/aes_core/SB1/n3184 ), .Y(\U1/aes_core/SB1/n3061 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB1/U1546  ( .A0(\U1/aes_core/SB1/n3185 ), 
        .A1(\U1/aes_core/SB1/n2968 ), .B0(\U1/aes_core/SB1/n3061 ), .B1(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n1733 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1545  ( .A0(\U1/aes_core/SB1/n3218 ), 
        .A1(\U1/aes_core/SB1/n3258 ), .B0(\U1/aes_core/SB1/n2983 ), .B1(
        \U1/aes_core/SB1/n3076 ), .C0(\U1/aes_core/SB1/n3220 ), .C1(
        \U1/aes_core/SB1/n3249 ), .Y(\U1/aes_core/SB1/n1732 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1544  ( .A(\U1/aes_core/SB1/n3079 ), .Y(
        \U1/aes_core/SB1/n3147 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1543  ( .A(\U1/aes_core/SB1/n3251 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3173 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1542  ( .A(\U1/aes_core/SB1/n3146 ), .B(
        \U1/aes_core/SB1/n2968 ), .Y(\U1/aes_core/SB1/n3000 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1541  ( .A(\U1/aes_core/SB1/n2982 ), .B(
        \U1/aes_core/SB1/n3189 ), .Y(\U1/aes_core/SB1/n3020 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1540  ( .A(\U1/aes_core/SB1/n3146 ), .B(
        \U1/aes_core/SB1/n3187 ), .Y(\U1/aes_core/SB1/n3119 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1539  ( .A(\U1/aes_core/SB1/n3173 ), .B(
        \U1/aes_core/SB1/n3000 ), .C(\U1/aes_core/SB1/n3020 ), .D(
        \U1/aes_core/SB1/n3119 ), .Y(\U1/aes_core/SB1/n1731 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1538  ( .A(\U1/aes_core/SB1/n3166 ), .B(
        \U1/aes_core/SB1/n3079 ), .Y(\U1/aes_core/SB1/n3042 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1537  ( .A(\U1/aes_core/SB1/n3152 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3052 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1536  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3068 ), .Y(\U1/aes_core/SB1/n3083 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1535  ( .AN(\U1/aes_core/SB1/n3042 ), 
        .B(\U1/aes_core/SB1/n3052 ), .C(\U1/aes_core/SB1/n3083 ), .Y(
        \U1/aes_core/SB1/n1730 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1534  ( .A(\U1/aes_core/SB1/n2977 ), .B(
        \U1/aes_core/SB1/n1734 ), .C(\U1/aes_core/SB1/n1733 ), .D(
        \U1/aes_core/SB1/n1732 ), .E(\U1/aes_core/SB1/n1731 ), .F(
        \U1/aes_core/SB1/n1730 ), .Y(\U1/aes_core/SB1/n3264 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1533  ( .A0(\U1/aes_core/SB1/n2982 ), 
        .A1(\U1/aes_core/SB1/n3210 ), .B0(\U1/aes_core/SB1/n3241 ), .Y(
        \U1/aes_core/SB1/n1735 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1532  ( .A(\U1/aes_core/SB1/n2968 ), .B(
        \U1/aes_core/SB1/n3068 ), .Y(\U1/aes_core/SB1/n3105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1531  ( .A(\U1/aes_core/SB1/n3185 ), .B(
        \U1/aes_core/SB1/n3233 ), .Y(\U1/aes_core/SB1/n2997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1530  ( .A(\U1/aes_core/SB1/n3233 ), .B(
        \U1/aes_core/SB1/n3189 ), .Y(\U1/aes_core/SB1/n3048 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1529  ( .A(\U1/aes_core/SB1/n1735 ), .B(
        \U1/aes_core/SB1/n3105 ), .C(\U1/aes_core/SB1/n2997 ), .D(
        \U1/aes_core/SB1/n3048 ), .Y(\U1/aes_core/SB1/n1739 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1528  ( .A0(\U1/aes_core/SB1/n3236 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n2983 ), .B1(
        \U1/aes_core/SB1/n3208 ), .C0(\U1/aes_core/SB1/n3237 ), .C1(
        \U1/aes_core/SB1/n3094 ), .Y(\U1/aes_core/SB1/n1738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1527  ( .A(\U1/aes_core/SB1/n3188 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n3029 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1526  ( .A(\U1/aes_core/SB1/n3187 ), .B(
        \U1/aes_core/SB1/n3239 ), .Y(\U1/aes_core/SB1/n3169 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1525  ( .A(\U1/aes_core/SB1/n3187 ), .B(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n3016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1524  ( .A(\U1/aes_core/SB1/n3242 ), .B(
        \U1/aes_core/SB1/n3232 ), .Y(\U1/aes_core/SB1/n2978 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1523  ( .A(\U1/aes_core/SB1/n3029 ), .B(
        \U1/aes_core/SB1/n3169 ), .C(\U1/aes_core/SB1/n3016 ), .D(
        \U1/aes_core/SB1/n2978 ), .Y(\U1/aes_core/SB1/n1737 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1522  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1521  ( .A(\U1/aes_core/SB1/n3251 ), .B(
        \U1/aes_core/SB1/n3212 ), .Y(\U1/aes_core/SB1/n3064 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1520  ( .A(\U1/aes_core/SB1/n3241 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1519  ( .A(\U1/aes_core/SB1/n2994 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n2965 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1518  ( .A(\U1/aes_core/SB1/n3091 ), .B(
        \U1/aes_core/SB1/n3064 ), .C(\U1/aes_core/SB1/n3115 ), .D(
        \U1/aes_core/SB1/n2965 ), .Y(\U1/aes_core/SB1/n1736 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1517  ( .A(\U1/aes_core/SB1/n1739 ), .B(
        \U1/aes_core/SB1/n1738 ), .C(\U1/aes_core/SB1/n1737 ), .D(
        \U1/aes_core/SB1/n1736 ), .Y(\U1/aes_core/SB1/n2892 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1516  ( .A(\U1/aes_core/SB1/n2346 ), .B(
        \U1/aes_core/SB1/n2903 ), .C(\U1/aes_core/SB1/n3264 ), .D(
        \U1/aes_core/SB1/n2892 ), .Y(\U1/aes_core/SB1/n1748 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1515  ( .A(\U1/aes_core/SB1/n3218 ), .Y(
        \U1/aes_core/SB1/n3142 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1514  ( .A0(\U1/aes_core/SB1/n3094 ), 
        .A1(\U1/aes_core/SB1/n2328 ), .B0(\U1/aes_core/SB1/n3063 ), .B1(
        \U1/aes_core/SB1/n3249 ), .Y(\U1/aes_core/SB1/n1740 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1513  ( .A0(\U1/aes_core/SB1/n3142 ), 
        .A1(\U1/aes_core/SB1/n3194 ), .B0(\U1/aes_core/SB1/n3243 ), .B1(
        \U1/aes_core/SB1/n3251 ), .C0(\U1/aes_core/SB1/n1740 ), .Y(
        \U1/aes_core/SB1/n1747 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1512  ( .A(\U1/aes_core/SB1/n3163 ), .B(
        \U1/aes_core/SB1/n3166 ), .Y(\U1/aes_core/SB1/n3162 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1511  ( .A0(\U1/aes_core/SB1/n3097 ), 
        .A1(\U1/aes_core/SB1/n3166 ), .B0(\U1/aes_core/SB1/n3079 ), .B1(
        \U1/aes_core/SB1/n3207 ), .Y(\U1/aes_core/SB1/n1741 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1510  ( .A0(\U1/aes_core/SB1/n2994 ), 
        .A1(\U1/aes_core/SB1/n3162 ), .B0(\U1/aes_core/SB1/n3213 ), .B1(
        \U1/aes_core/SB1/n3232 ), .C0(\U1/aes_core/SB1/n1741 ), .Y(
        \U1/aes_core/SB1/n1746 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1509  ( .A(\U1/aes_core/SB1/n3237 ), .B(
        \U1/aes_core/SB1/n3096 ), .Y(\U1/aes_core/SB1/n1744 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1508  ( .A(\U1/aes_core/SB1/n3187 ), .B(
        \U1/aes_core/SB1/n3212 ), .Y(\U1/aes_core/SB1/n3154 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1507  ( .A(\U1/aes_core/SB1/n3154 ), .Y(
        \U1/aes_core/SB1/n1743 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1506  ( .A(\U1/aes_core/SB1/n3145 ), .B(
        \U1/aes_core/SB1/n3218 ), .Y(\U1/aes_core/SB1/n3026 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1505  ( .A(\U1/aes_core/SB1/n3223 ), .B(
        \U1/aes_core/SB1/n3221 ), .Y(\U1/aes_core/SB1/n3179 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1503  ( .A(\U1/aes_core/SB1/n3194 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3036 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1501  ( .A0(\U1/aes_core/SB1/n3153 ), 
        .A1(\U1/aes_core/SB1/n1744 ), .B0(\U1/aes_core/SB1/n3130 ), .B1(
        \U1/aes_core/SB1/n1743 ), .C0(\U1/aes_core/SB1/n1742 ), .Y(
        \U1/aes_core/SB1/n1745 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1500  ( .AN(\U1/aes_core/SB1/n1748 ), 
        .B(\U1/aes_core/SB1/n1747 ), .C(\U1/aes_core/SB1/n1746 ), .D(
        \U1/aes_core/SB1/n1745 ), .Y(\U1/aes_core/sb1 [0]) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1499  ( .A(Dout[78]), .Y(
        \U1/aes_core/SB1/n1755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1498  ( .A(Dout[79]), .Y(
        \U1/aes_core/SB1/n1750 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1497  ( .A(\U1/aes_core/SB1/n1755 ), .B(
        \U1/aes_core/SB1/n1750 ), .Y(\U1/aes_core/SB1/n1760 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1496  ( .A(Dout[77]), .Y(
        \U1/aes_core/SB1/n1749 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1495  ( .A(\U1/aes_core/SB1/n1749 ), .B(
        Dout[76]), .Y(\U1/aes_core/SB1/n1767 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1494  ( .A(\U1/aes_core/SB1/n1760 ), .B(
        \U1/aes_core/SB1/n1767 ), .Y(\U1/aes_core/SB1/n3300 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1493  ( .A(Dout[75]), .Y(
        \U1/aes_core/SB1/n1758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1492  ( .A(\U1/aes_core/SB1/n1758 ), .B(
        Dout[74]), .Y(\U1/aes_core/SB1/n1773 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1491  ( .A(Dout[72]), .Y(
        \U1/aes_core/SB1/n1751 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1490  ( .A(\U1/aes_core/SB1/n1751 ), .B(
        Dout[73]), .Y(\U1/aes_core/SB1/n1761 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1489  ( .A(\U1/aes_core/SB1/n1773 ), .B(
        \U1/aes_core/SB1/n1761 ), .Y(\U1/aes_core/SB1/n1912 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1488  ( .A(\U1/aes_core/SB1/n3300 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n1821 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1487  ( .A(Dout[73]), .Y(
        \U1/aes_core/SB1/n1752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1486  ( .A(\U1/aes_core/SB1/n1752 ), .B(
        Dout[72]), .Y(\U1/aes_core/SB1/n1770 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1485  ( .A(Dout[74]), .Y(
        \U1/aes_core/SB1/n1757 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1484  ( .A(\U1/aes_core/SB1/n1757 ), .B(
        Dout[75]), .Y(\U1/aes_core/SB1/n1754 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1483  ( .A(\U1/aes_core/SB1/n1770 ), .B(
        \U1/aes_core/SB1/n1754 ), .Y(\U1/aes_core/SB1/n3346 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1482  ( .A(Dout[76]), .Y(
        \U1/aes_core/SB1/n1753 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1481  ( .A(\U1/aes_core/SB1/n1749 ), .B(
        \U1/aes_core/SB1/n1753 ), .Y(\U1/aes_core/SB1/n1781 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1480  ( .A(\U1/aes_core/SB1/n1750 ), .B(
        Dout[78]), .Y(\U1/aes_core/SB1/n1756 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1479  ( .A(\U1/aes_core/SB1/n1781 ), .B(
        \U1/aes_core/SB1/n1756 ), .Y(\U1/aes_core/SB1/n2021 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1478  ( .A0(\U1/aes_core/SB1/n1912 ), 
        .A1(\U1/aes_core/SB1/n3346 ), .B0(\U1/aes_core/SB1/n2021 ), .Y(
        \U1/aes_core/SB1/n1766 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1477  ( .A(\U1/aes_core/SB1/n1752 ), .B(
        \U1/aes_core/SB1/n1751 ), .Y(\U1/aes_core/SB1/n1772 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1476  ( .A(\U1/aes_core/SB1/n1754 ), .B(
        \U1/aes_core/SB1/n1772 ), .Y(\U1/aes_core/SB1/n2020 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1475  ( .A(\U1/aes_core/SB1/n1753 ), .B(
        Dout[77]), .Y(\U1/aes_core/SB1/n1783 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1474  ( .A(\U1/aes_core/SB1/n1760 ), .B(
        \U1/aes_core/SB1/n1783 ), .Y(\U1/aes_core/SB1/n1995 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1473  ( .A(Dout[75]), .B(Dout[74]), .Y(
        \U1/aes_core/SB1/n1780 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1472  ( .A(\U1/aes_core/SB1/n1772 ), .B(
        \U1/aes_core/SB1/n1780 ), .Y(\U1/aes_core/SB1/n3301 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1471  ( .A(\U1/aes_core/SB1/n3301 ), .Y(
        \U1/aes_core/SB1/n3339 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1470  ( .A(Dout[73]), .B(Dout[72]), .Y(
        \U1/aes_core/SB1/n1779 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1469  ( .A(\U1/aes_core/SB1/n1754 ), .B(
        \U1/aes_core/SB1/n1779 ), .Y(\U1/aes_core/SB1/n3296 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1468  ( .A(\U1/aes_core/SB1/n3296 ), .Y(
        \U1/aes_core/SB1/n3333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1467  ( .A(\U1/aes_core/SB1/n3339 ), .B(
        \U1/aes_core/SB1/n3333 ), .Y(\U1/aes_core/SB1/n1823 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1466  ( .A(Dout[79]), .B(Dout[78]), .Y(
        \U1/aes_core/SB1/n1774 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1465  ( .A(\U1/aes_core/SB1/n1767 ), .B(
        \U1/aes_core/SB1/n1774 ), .Y(\U1/aes_core/SB1/n3309 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1464  ( .A0(\U1/aes_core/SB1/n2020 ), 
        .A1(\U1/aes_core/SB1/n1995 ), .B0(\U1/aes_core/SB1/n1823 ), .B1(
        \U1/aes_core/SB1/n3309 ), .Y(\U1/aes_core/SB1/n1765 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1463  ( .A(\U1/aes_core/SB1/n1754 ), .B(
        \U1/aes_core/SB1/n1761 ), .Y(\U1/aes_core/SB1/n1888 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1462  ( .A(\U1/aes_core/SB1/n1767 ), .B(
        \U1/aes_core/SB1/n1756 ), .Y(\U1/aes_core/SB1/n3344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1461  ( .A(Dout[77]), .B(Dout[76]), .Y(
        \U1/aes_core/SB1/n1759 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1460  ( .A(\U1/aes_core/SB1/n1760 ), .B(
        \U1/aes_core/SB1/n1759 ), .Y(\U1/aes_core/SB1/n3280 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1459  ( .A(\U1/aes_core/SB1/n1783 ), .B(
        \U1/aes_core/SB1/n1756 ), .Y(\U1/aes_core/SB1/n3278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1458  ( .A(\U1/aes_core/SB1/n1773 ), .B(
        \U1/aes_core/SB1/n1779 ), .Y(\U1/aes_core/SB1/n2010 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1457  ( .A0(\U1/aes_core/SB1/n1888 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n3301 ), .B1(
        \U1/aes_core/SB1/n3280 ), .C0(\U1/aes_core/SB1/n3278 ), .C1(
        \U1/aes_core/SB1/n2010 ), .Y(\U1/aes_core/SB1/n1764 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1456  ( .A(\U1/aes_core/SB1/n1755 ), .B(
        Dout[79]), .Y(\U1/aes_core/SB1/n1782 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1455  ( .A(\U1/aes_core/SB1/n1782 ), .B(
        \U1/aes_core/SB1/n1759 ), .Y(\U1/aes_core/SB1/n3308 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1454  ( .A(\U1/aes_core/SB1/n3308 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n1873 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1453  ( .A(\U1/aes_core/SB1/n1770 ), .B(
        \U1/aes_core/SB1/n1773 ), .Y(\U1/aes_core/SB1/n3342 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1452  ( .A(\U1/aes_core/SB1/n3342 ), .Y(
        \U1/aes_core/SB1/n2058 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1451  ( .A(\U1/aes_core/SB1/n1759 ), .B(
        \U1/aes_core/SB1/n1756 ), .Y(\U1/aes_core/SB1/n1806 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1450  ( .A(\U1/aes_core/SB1/n1806 ), .Y(
        \U1/aes_core/SB1/n3268 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1449  ( .A(\U1/aes_core/SB1/n2058 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n1856 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1448  ( .A(\U1/aes_core/SB1/n1758 ), .B(
        \U1/aes_core/SB1/n1757 ), .Y(\U1/aes_core/SB1/n1769 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1447  ( .A(\U1/aes_core/SB1/n1772 ), .B(
        \U1/aes_core/SB1/n1769 ), .Y(\U1/aes_core/SB1/n2006 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1446  ( .A(\U1/aes_core/SB1/n2006 ), .Y(
        \U1/aes_core/SB1/n2068 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U1445  ( .A(\U1/aes_core/SB1/n1774 ), .B(
        \U1/aes_core/SB1/n1759 ), .Y(\U1/aes_core/SB1/n3299 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1444  ( .A(\U1/aes_core/SB1/n2068 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1928 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1443  ( .A(\U1/aes_core/SB1/n1760 ), .B(
        \U1/aes_core/SB1/n1781 ), .Y(\U1/aes_core/SB1/n3347 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1442  ( .A(\U1/aes_core/SB1/n3347 ), .Y(
        \U1/aes_core/SB1/n3305 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1441  ( .A(\U1/aes_core/SB1/n3305 ), .B(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n1953 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1440  ( .AN(\U1/aes_core/SB1/n1873 ), 
        .B(\U1/aes_core/SB1/n1856 ), .C(\U1/aes_core/SB1/n1928 ), .D(
        \U1/aes_core/SB1/n1953 ), .Y(\U1/aes_core/SB1/n1763 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1439  ( .A(\U1/aes_core/SB1/n1995 ), .Y(
        \U1/aes_core/SB1/n3269 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1438  ( .A(\U1/aes_core/SB1/n1780 ), .B(
        \U1/aes_core/SB1/n1761 ), .Y(\U1/aes_core/SB1/n2017 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1437  ( .A(\U1/aes_core/SB1/n2017 ), .Y(
        \U1/aes_core/SB1/n2054 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1436  ( .A(\U1/aes_core/SB1/n3269 ), .B(
        \U1/aes_core/SB1/n2054 ), .Y(\U1/aes_core/SB1/n1843 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1435  ( .A(\U1/aes_core/SB1/n3278 ), .Y(
        \U1/aes_core/SB1/n3332 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1434  ( .A(\U1/aes_core/SB1/n1761 ), .B(
        \U1/aes_core/SB1/n1769 ), .Y(\U1/aes_core/SB1/n2057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1433  ( .A(\U1/aes_core/SB1/n2057 ), .Y(
        \U1/aes_core/SB1/n2019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1432  ( .A(\U1/aes_core/SB1/n3332 ), .B(
        \U1/aes_core/SB1/n2019 ), .Y(\U1/aes_core/SB1/n1879 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1431  ( .A(\U1/aes_core/SB1/n3269 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1966 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U1430  ( .A(\U1/aes_core/SB1/n1843 ), .B(
        \U1/aes_core/SB1/n1879 ), .C(\U1/aes_core/SB1/n1966 ), .Y(
        \U1/aes_core/SB1/n1762 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1429  ( .A(\U1/aes_core/SB1/n1821 ), .B(
        \U1/aes_core/SB1/n1766 ), .C(\U1/aes_core/SB1/n1765 ), .D(
        \U1/aes_core/SB1/n1764 ), .E(\U1/aes_core/SB1/n1763 ), .F(
        \U1/aes_core/SB1/n1762 ), .Y(\U1/aes_core/SB1/n3353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1428  ( .A(\U1/aes_core/SB1/n1995 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n1944 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1427  ( .A(\U1/aes_core/SB1/n2010 ), .Y(
        \U1/aes_core/SB1/n3330 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1426  ( .A(\U1/aes_core/SB1/n1888 ), .Y(
        \U1/aes_core/SB1/n3334 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1425  ( .A(\U1/aes_core/SB1/n1767 ), .B(
        \U1/aes_core/SB1/n1782 ), .Y(\U1/aes_core/SB1/n3343 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1424  ( .A(\U1/aes_core/SB1/n3343 ), .Y(
        \U1/aes_core/SB1/n3274 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1423  ( .A0(\U1/aes_core/SB1/n3330 ), 
        .A1(\U1/aes_core/SB1/n3334 ), .B0(\U1/aes_core/SB1/n3274 ), .Y(
        \U1/aes_core/SB1/n1768 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1422  ( .A(\U1/aes_core/SB1/n3305 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1903 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1421  ( .A(\U1/aes_core/SB1/n2021 ), .Y(
        \U1/aes_core/SB1/n2053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1420  ( .A(\U1/aes_core/SB1/n3339 ), .B(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n1865 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1419  ( .AN(\U1/aes_core/SB1/n1944 ), 
        .B(\U1/aes_core/SB1/n1768 ), .C(\U1/aes_core/SB1/n1903 ), .D(
        \U1/aes_core/SB1/n1865 ), .Y(\U1/aes_core/SB1/n1778 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1418  ( .A(\U1/aes_core/SB1/n3309 ), .Y(
        \U1/aes_core/SB1/n1976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1417  ( .A(\U1/aes_core/SB1/n1770 ), .B(
        \U1/aes_core/SB1/n1780 ), .Y(\U1/aes_core/SB1/n2039 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1416  ( .A(\U1/aes_core/SB1/n2039 ), .Y(
        \U1/aes_core/SB1/n3340 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1415  ( .A(\U1/aes_core/SB1/n3280 ), .Y(
        \U1/aes_core/SB1/n2055 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1414  ( .A(\U1/aes_core/SB1/n1779 ), .B(
        \U1/aes_core/SB1/n1769 ), .Y(\U1/aes_core/SB1/n3281 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1413  ( .A(\U1/aes_core/SB1/n3281 ), .Y(
        \U1/aes_core/SB1/n3331 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U1412  ( .A0(\U1/aes_core/SB1/n1976 ), 
        .A1(\U1/aes_core/SB1/n2068 ), .B0(\U1/aes_core/SB1/n3340 ), .B1(
        \U1/aes_core/SB1/n2055 ), .C0(\U1/aes_core/SB1/n3331 ), .C1(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n1777 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1411  ( .A(\U1/aes_core/SB1/n3300 ), .Y(
        \U1/aes_core/SB1/n1952 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1410  ( .A(\U1/aes_core/SB1/n1774 ), .B(
        \U1/aes_core/SB1/n1781 ), .Y(\U1/aes_core/SB1/n2070 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1409  ( .A(\U1/aes_core/SB1/n1770 ), .B(
        \U1/aes_core/SB1/n1769 ), .Y(\U1/aes_core/SB1/n3279 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1408  ( .A0(\U1/aes_core/SB1/n2070 ), 
        .A1(\U1/aes_core/SB1/n3346 ), .B0(\U1/aes_core/SB1/n3279 ), .B1(
        \U1/aes_core/SB1/n1995 ), .Y(\U1/aes_core/SB1/n1771 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1407  ( .A0(\U1/aes_core/SB1/n2058 ), 
        .A1(\U1/aes_core/SB1/n3305 ), .B0(\U1/aes_core/SB1/n1952 ), .B1(
        \U1/aes_core/SB1/n2019 ), .C0(\U1/aes_core/SB1/n1771 ), .Y(
        \U1/aes_core/SB1/n1776 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1406  ( .A(\U1/aes_core/SB1/n3268 ), .B(
        \U1/aes_core/SB1/n2019 ), .Y(\U1/aes_core/SB1/n1880 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1405  ( .A(\U1/aes_core/SB1/n1773 ), .B(
        \U1/aes_core/SB1/n1772 ), .Y(\U1/aes_core/SB1/n3302 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1404  ( .A(\U1/aes_core/SB1/n3302 ), .Y(
        \U1/aes_core/SB1/n3276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1403  ( .A(\U1/aes_core/SB1/n3276 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n1845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1402  ( .A(\U1/aes_core/SB1/n2070 ), .Y(
        \U1/aes_core/SB1/n3324 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1401  ( .A(\U1/aes_core/SB1/n3324 ), .B(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n1929 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1400  ( .A(\U1/aes_core/SB1/n1783 ), .B(
        \U1/aes_core/SB1/n1774 ), .Y(\U1/aes_core/SB1/n2065 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1399  ( .A(\U1/aes_core/SB1/n2065 ), .Y(
        \U1/aes_core/SB1/n3322 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1398  ( .A(\U1/aes_core/SB1/n3322 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1852 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB1/U1397  ( .A(\U1/aes_core/SB1/n1880 ), .B(
        \U1/aes_core/SB1/n1845 ), .C(\U1/aes_core/SB1/n1929 ), .D(
        \U1/aes_core/SB1/n1852 ), .Y(\U1/aes_core/SB1/n1775 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1396  ( .AN(\U1/aes_core/SB1/n1778 ), 
        .B(\U1/aes_core/SB1/n1777 ), .C(\U1/aes_core/SB1/n1776 ), .D(
        \U1/aes_core/SB1/n1775 ), .Y(\U1/aes_core/SB1/n3295 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1395  ( .A(\U1/aes_core/SB1/n1780 ), .B(
        \U1/aes_core/SB1/n1779 ), .Y(\U1/aes_core/SB1/n3297 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1394  ( .A(\U1/aes_core/SB1/n3297 ), .B(
        \U1/aes_core/SB1/n2021 ), .Y(\U1/aes_core/SB1/n1965 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1393  ( .A(\U1/aes_core/SB1/n3300 ), .B(
        \U1/aes_core/SB1/n2006 ), .Y(\U1/aes_core/SB1/n1878 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1392  ( .A(\U1/aes_core/SB1/n3333 ), .B(
        \U1/aes_core/SB1/n3305 ), .Y(\U1/aes_core/SB1/n1842 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1391  ( .A0(\U1/aes_core/SB1/n3300 ), 
        .A1(\U1/aes_core/SB1/n3342 ), .B0(\U1/aes_core/SB1/n1842 ), .Y(
        \U1/aes_core/SB1/n1787 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1390  ( .A(\U1/aes_core/SB1/n1912 ), .Y(
        \U1/aes_core/SB1/n3325 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1389  ( .A(\U1/aes_core/SB1/n3268 ), .B(
        \U1/aes_core/SB1/n3325 ), .Y(\U1/aes_core/SB1/n1977 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1388  ( .A(\U1/aes_core/SB1/n3268 ), .B(
        \U1/aes_core/SB1/n3334 ), .Y(\U1/aes_core/SB1/n1954 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1387  ( .A(\U1/aes_core/SB1/n1782 ), .B(
        \U1/aes_core/SB1/n1781 ), .Y(\U1/aes_core/SB1/n2008 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1386  ( .A(\U1/aes_core/SB1/n2008 ), .Y(
        \U1/aes_core/SB1/n3307 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1385  ( .A(\U1/aes_core/SB1/n3307 ), .B(
        \U1/aes_core/SB1/n2019 ), .Y(\U1/aes_core/SB1/n1855 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1384  ( .A(\U1/aes_core/SB1/n3307 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1902 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1383  ( .A(\U1/aes_core/SB1/n1977 ), .B(
        \U1/aes_core/SB1/n1954 ), .C(\U1/aes_core/SB1/n1855 ), .D(
        \U1/aes_core/SB1/n1902 ), .Y(\U1/aes_core/SB1/n1786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1382  ( .A(\U1/aes_core/SB1/n3346 ), .Y(
        \U1/aes_core/SB1/n3275 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1381  ( .A(\U1/aes_core/SB1/n3275 ), .B(
        \U1/aes_core/SB1/n1976 ), .Y(\U1/aes_core/SB1/n1927 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1380  ( .A(\U1/aes_core/SB1/n3297 ), .Y(
        \U1/aes_core/SB1/n3282 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1379  ( .A(\U1/aes_core/SB1/n1976 ), .B(
        \U1/aes_core/SB1/n3282 ), .Y(\U1/aes_core/SB1/n1922 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1378  ( .A(\U1/aes_core/SB1/n3322 ), .B(
        \U1/aes_core/SB1/n3276 ), .Y(\U1/aes_core/SB1/n1830 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1377  ( .A(\U1/aes_core/SB1/n3299 ), .B(
        \U1/aes_core/SB1/n2019 ), .Y(\U1/aes_core/SB1/n1909 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1376  ( .A(\U1/aes_core/SB1/n1927 ), .B(
        \U1/aes_core/SB1/n1922 ), .C(\U1/aes_core/SB1/n1830 ), .D(
        \U1/aes_core/SB1/n1909 ), .Y(\U1/aes_core/SB1/n1785 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1375  ( .A(\U1/aes_core/SB1/n3279 ), .Y(
        \U1/aes_core/SB1/n3323 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1374  ( .A(\U1/aes_core/SB1/n3274 ), .B(
        \U1/aes_core/SB1/n3323 ), .Y(\U1/aes_core/SB1/n1820 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1373  ( .A(\U1/aes_core/SB1/n2054 ), .B(
        \U1/aes_core/SB1/n3274 ), .Y(\U1/aes_core/SB1/n1864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1372  ( .A(\U1/aes_core/SB1/n1783 ), .B(
        \U1/aes_core/SB1/n1782 ), .Y(\U1/aes_core/SB1/n3303 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1371  ( .A(\U1/aes_core/SB1/n3303 ), .Y(
        \U1/aes_core/SB1/n3329 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1370  ( .A(\U1/aes_core/SB1/n2068 ), .B(
        \U1/aes_core/SB1/n3329 ), .Y(\U1/aes_core/SB1/n1890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1369  ( .A(\U1/aes_core/SB1/n2054 ), .B(
        \U1/aes_core/SB1/n3324 ), .Y(\U1/aes_core/SB1/n1990 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1368  ( .A(\U1/aes_core/SB1/n1820 ), .B(
        \U1/aes_core/SB1/n1864 ), .C(\U1/aes_core/SB1/n1890 ), .D(
        \U1/aes_core/SB1/n1990 ), .Y(\U1/aes_core/SB1/n1784 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1367  ( .A(\U1/aes_core/SB1/n1965 ), .B(
        \U1/aes_core/SB1/n1878 ), .C(\U1/aes_core/SB1/n1787 ), .D(
        \U1/aes_core/SB1/n1786 ), .E(\U1/aes_core/SB1/n1785 ), .F(
        \U1/aes_core/SB1/n1784 ), .Y(\U1/aes_core/SB1/n3286 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1366  ( .A(\U1/aes_core/SB1/n3279 ), .B(
        \U1/aes_core/SB1/n2021 ), .Y(\U1/aes_core/SB1/n1831 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1365  ( .A(\U1/aes_core/SB1/n3280 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n1980 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1364  ( .A(\U1/aes_core/SB1/n3278 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n1872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1363  ( .A(\U1/aes_core/SB1/n3278 ), .B(
        \U1/aes_core/SB1/n3281 ), .Y(\U1/aes_core/SB1/n1881 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1362  ( .A(\U1/aes_core/SB1/n3342 ), .B(
        \U1/aes_core/SB1/n3308 ), .Y(\U1/aes_core/SB1/n1919 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1361  ( .A(\U1/aes_core/SB1/n3307 ), .B(
        \U1/aes_core/SB1/n3325 ), .Y(\U1/aes_core/SB1/n1923 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1360  ( .A(\U1/aes_core/SB1/n2058 ), .B(
        \U1/aes_core/SB1/n3329 ), .Y(\U1/aes_core/SB1/n1844 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1359  ( .A(\U1/aes_core/SB1/n3331 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1857 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1358  ( .AN(\U1/aes_core/SB1/n1919 ), 
        .B(\U1/aes_core/SB1/n1923 ), .C(\U1/aes_core/SB1/n1844 ), .D(
        \U1/aes_core/SB1/n1857 ), .Y(\U1/aes_core/SB1/n1791 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1357  ( .A(\U1/aes_core/SB1/n3300 ), .B(
        \U1/aes_core/SB1/n3281 ), .Y(\U1/aes_core/SB1/n1891 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1356  ( .A(\U1/aes_core/SB1/n3347 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n1967 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1355  ( .A(\U1/aes_core/SB1/n1995 ), .B(
        \U1/aes_core/SB1/n3346 ), .Y(\U1/aes_core/SB1/n1930 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1354  ( .A(\U1/aes_core/SB1/n1995 ), .B(
        \U1/aes_core/SB1/n2006 ), .Y(\U1/aes_core/SB1/n1828 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1353  ( .A0(\U1/aes_core/SB1/n3281 ), 
        .A1(\U1/aes_core/SB1/n1995 ), .B0(\U1/aes_core/SB1/n3300 ), .B1(
        \U1/aes_core/SB1/n3346 ), .Y(\U1/aes_core/SB1/n1789 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1352  ( .A0(\U1/aes_core/SB1/n1888 ), 
        .A1(\U1/aes_core/SB1/n2070 ), .B0(\U1/aes_core/SB1/n2020 ), .B1(
        \U1/aes_core/SB1/n3280 ), .Y(\U1/aes_core/SB1/n1788 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1351  ( .A(\U1/aes_core/SB1/n1891 ), .B(
        \U1/aes_core/SB1/n1967 ), .C(\U1/aes_core/SB1/n1930 ), .D(
        \U1/aes_core/SB1/n1828 ), .E(\U1/aes_core/SB1/n1789 ), .F(
        \U1/aes_core/SB1/n1788 ), .Y(\U1/aes_core/SB1/n1790 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1350  ( .A(\U1/aes_core/SB1/n1831 ), .B(
        \U1/aes_core/SB1/n1980 ), .C(\U1/aes_core/SB1/n1872 ), .D(
        \U1/aes_core/SB1/n1881 ), .E(\U1/aes_core/SB1/n1791 ), .F(
        \U1/aes_core/SB1/n1790 ), .Y(\U1/aes_core/SB1/n3321 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U1349  ( .A1N(\U1/aes_core/SB1/n3299 ), 
        .A0(\U1/aes_core/SB1/n3343 ), .B0(\U1/aes_core/SB1/n2020 ), .Y(
        \U1/aes_core/SB1/n1792 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1348  ( .A(\U1/aes_core/SB1/n1995 ), .B(
        \U1/aes_core/SB1/n2039 ), .Y(\U1/aes_core/SB1/n1943 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1347  ( .A(\U1/aes_core/SB1/n3280 ), .B(
        \U1/aes_core/SB1/n2057 ), .Y(\U1/aes_core/SB1/n1850 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1346  ( .A(\U1/aes_core/SB1/n3280 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n1886 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1345  ( .A(\U1/aes_core/SB1/n1792 ), .B(
        \U1/aes_core/SB1/n1943 ), .C(\U1/aes_core/SB1/n1850 ), .D(
        \U1/aes_core/SB1/n1886 ), .Y(\U1/aes_core/SB1/n1797 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1344  ( .A0(\U1/aes_core/SB1/n2057 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n2021 ), .B1(
        \U1/aes_core/SB1/n3296 ), .C0(\U1/aes_core/SB1/n1912 ), .C1(
        \U1/aes_core/SB1/n3309 ), .Y(\U1/aes_core/SB1/n1796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1343  ( .A(\U1/aes_core/SB1/n3342 ), .B(
        \U1/aes_core/SB1/n3309 ), .Y(\U1/aes_core/SB1/n1972 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1342  ( .A(\U1/aes_core/SB1/n2065 ), .B(
        \U1/aes_core/SB1/n2010 ), .Y(\U1/aes_core/SB1/n1833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1341  ( .A(\U1/aes_core/SB1/n1833 ), .Y(
        \U1/aes_core/SB1/n1793 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1340  ( .A(\U1/aes_core/SB1/n3329 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1339  ( .A(\U1/aes_core/SB1/n1976 ), .B(
        \U1/aes_core/SB1/n2054 ), .Y(\U1/aes_core/SB1/n1853 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1338  ( .AN(\U1/aes_core/SB1/n1972 ), 
        .B(\U1/aes_core/SB1/n1793 ), .C(\U1/aes_core/SB1/n1866 ), .D(
        \U1/aes_core/SB1/n1853 ), .Y(\U1/aes_core/SB1/n1795 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1337  ( .A(\U1/aes_core/SB1/n1888 ), .B(
        \U1/aes_core/SB1/n2021 ), .Y(\U1/aes_core/SB1/n1918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1336  ( .A(\U1/aes_core/SB1/n1806 ), .B(
        \U1/aes_core/SB1/n3297 ), .Y(\U1/aes_core/SB1/n1895 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1335  ( .A(\U1/aes_core/SB1/n2008 ), .B(
        \U1/aes_core/SB1/n2020 ), .Y(\U1/aes_core/SB1/n1935 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1334  ( .A(\U1/aes_core/SB1/n2008 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n1827 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1333  ( .A(\U1/aes_core/SB1/n1918 ), .B(
        \U1/aes_core/SB1/n1895 ), .C(\U1/aes_core/SB1/n1935 ), .D(
        \U1/aes_core/SB1/n1827 ), .Y(\U1/aes_core/SB1/n1794 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1332  ( .A(\U1/aes_core/SB1/n1797 ), .B(
        \U1/aes_core/SB1/n1796 ), .C(\U1/aes_core/SB1/n1795 ), .D(
        \U1/aes_core/SB1/n1794 ), .Y(\U1/aes_core/SB1/n3293 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1331  ( .A(\U1/aes_core/SB1/n3308 ), .Y(
        \U1/aes_core/SB1/n3327 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1330  ( .A0(\U1/aes_core/SB1/n3330 ), 
        .A1(\U1/aes_core/SB1/n3268 ), .B0(\U1/aes_core/SB1/n2068 ), .B1(
        \U1/aes_core/SB1/n3327 ), .Y(\U1/aes_core/SB1/n1798 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1329  ( .A0(\U1/aes_core/SB1/n3297 ), 
        .A1(\U1/aes_core/SB1/n3347 ), .B0(\U1/aes_core/SB1/n3280 ), .B1(
        \U1/aes_core/SB1/n3346 ), .C0(\U1/aes_core/SB1/n1798 ), .Y(
        \U1/aes_core/SB1/n1804 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1328  ( .A(\U1/aes_core/SB1/n3303 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n1862 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1327  ( .A(\U1/aes_core/SB1/n3332 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1326  ( .A(\U1/aes_core/SB1/n3268 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1325  ( .A(\U1/aes_core/SB1/n3330 ), .B(
        \U1/aes_core/SB1/n3307 ), .Y(\U1/aes_core/SB1/n1839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1324  ( .AN(\U1/aes_core/SB1/n1862 ), 
        .B(\U1/aes_core/SB1/n1874 ), .C(\U1/aes_core/SB1/n1867 ), .D(
        \U1/aes_core/SB1/n1839 ), .Y(\U1/aes_core/SB1/n1803 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1323  ( .A(\U1/aes_core/SB1/n3281 ), .B(
        \U1/aes_core/SB1/n2057 ), .Y(\U1/aes_core/SB1/n1948 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1322  ( .A0(\U1/aes_core/SB1/n3325 ), 
        .A1(\U1/aes_core/SB1/n1948 ), .B0(\U1/aes_core/SB1/n3322 ), .Y(
        \U1/aes_core/SB1/n1801 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1321  ( .A(\U1/aes_core/SB1/n3344 ), .Y(
        \U1/aes_core/SB1/n1949 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1320  ( .A0(\U1/aes_core/SB1/n2058 ), 
        .A1(\U1/aes_core/SB1/n3323 ), .B0(\U1/aes_core/SB1/n1949 ), .Y(
        \U1/aes_core/SB1/n1800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1319  ( .A(\U1/aes_core/SB1/n2020 ), .Y(
        \U1/aes_core/SB1/n2060 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1318  ( .A0(\U1/aes_core/SB1/n1952 ), 
        .A1(\U1/aes_core/SB1/n1976 ), .B0(\U1/aes_core/SB1/n2060 ), .Y(
        \U1/aes_core/SB1/n1799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1317  ( .A(\U1/aes_core/SB1/n2058 ), .B(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n1925 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1316  ( .A(\U1/aes_core/SB1/n1801 ), .B(
        \U1/aes_core/SB1/n1800 ), .C(\U1/aes_core/SB1/n1799 ), .D(
        \U1/aes_core/SB1/n1925 ), .Y(\U1/aes_core/SB1/n1802 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1315  ( .A(\U1/aes_core/SB1/n3286 ), .B(
        \U1/aes_core/SB1/n3321 ), .C(\U1/aes_core/SB1/n3293 ), .D(
        \U1/aes_core/SB1/n1804 ), .E(\U1/aes_core/SB1/n1803 ), .F(
        \U1/aes_core/SB1/n1802 ), .Y(\U1/aes_core/SB1/n2074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1314  ( .A0(\U1/aes_core/SB1/n2019 ), 
        .A1(\U1/aes_core/SB1/n3330 ), .B0(\U1/aes_core/SB1/n3324 ), .Y(
        \U1/aes_core/SB1/n1805 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1313  ( .A(\U1/aes_core/SB1/n3269 ), .B(
        \U1/aes_core/SB1/n2058 ), .Y(\U1/aes_core/SB1/n1910 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1312  ( .A(\U1/aes_core/SB1/n2055 ), .B(
        \U1/aes_core/SB1/n3276 ), .Y(\U1/aes_core/SB1/n1819 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1311  ( .A(\U1/aes_core/SB1/n3340 ), .B(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n1921 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1310  ( .A(\U1/aes_core/SB1/n1805 ), .B(
        \U1/aes_core/SB1/n1910 ), .C(\U1/aes_core/SB1/n1819 ), .D(
        \U1/aes_core/SB1/n1921 ), .Y(\U1/aes_core/SB1/n1810 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1309  ( .A0(\U1/aes_core/SB1/n2020 ), 
        .A1(\U1/aes_core/SB1/n1806 ), .B0(\U1/aes_core/SB1/n3302 ), .B1(
        \U1/aes_core/SB1/n3347 ), .C0(\U1/aes_core/SB1/n3346 ), .C1(
        \U1/aes_core/SB1/n2065 ), .Y(\U1/aes_core/SB1/n1809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1308  ( .A(\U1/aes_core/SB1/n1976 ), .B(
        \U1/aes_core/SB1/n3334 ), .Y(\U1/aes_core/SB1/n1841 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1307  ( .A(\U1/aes_core/SB1/n2058 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1964 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1306  ( .A(\U1/aes_core/SB1/n3275 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1863 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1305  ( .A(\U1/aes_core/SB1/n3340 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1926 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1304  ( .A(\U1/aes_core/SB1/n1841 ), .B(
        \U1/aes_core/SB1/n1964 ), .C(\U1/aes_core/SB1/n1863 ), .D(
        \U1/aes_core/SB1/n1926 ), .Y(\U1/aes_core/SB1/n1808 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1303  ( .A(\U1/aes_core/SB1/n3340 ), .B(
        \U1/aes_core/SB1/n3332 ), .Y(\U1/aes_core/SB1/n1889 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1302  ( .A(\U1/aes_core/SB1/n3333 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n1876 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1301  ( .A(\U1/aes_core/SB1/n3274 ), .B(
        \U1/aes_core/SB1/n3276 ), .Y(\U1/aes_core/SB1/n1854 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1300  ( .A(\U1/aes_core/SB1/n3323 ), .B(
        \U1/aes_core/SB1/n3327 ), .Y(\U1/aes_core/SB1/n1829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1299  ( .A(\U1/aes_core/SB1/n1889 ), .B(
        \U1/aes_core/SB1/n1876 ), .C(\U1/aes_core/SB1/n1854 ), .D(
        \U1/aes_core/SB1/n1829 ), .Y(\U1/aes_core/SB1/n1807 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1298  ( .A(\U1/aes_core/SB1/n1810 ), .B(
        \U1/aes_core/SB1/n1809 ), .C(\U1/aes_core/SB1/n1808 ), .D(
        \U1/aes_core/SB1/n1807 ), .Y(\U1/aes_core/SB1/n1811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1297  ( .A(\U1/aes_core/SB1/n1811 ), .Y(
        \U1/aes_core/SB1/n3284 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1296  ( .A0(\U1/aes_core/SB1/n3308 ), 
        .A1(\U1/aes_core/SB1/n2039 ), .B0(\U1/aes_core/SB1/n3297 ), .B1(
        \U1/aes_core/SB1/n2070 ), .C0(\U1/aes_core/SB1/n3284 ), .Y(
        \U1/aes_core/SB1/n1818 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1295  ( .A(\U1/aes_core/SB1/n3329 ), .B(
        \U1/aes_core/SB1/n3274 ), .Y(\U1/aes_core/SB1/n1920 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U1294  ( .A1N(\U1/aes_core/SB1/n1920 ), 
        .A0(\U1/aes_core/SB1/n3305 ), .B0(\U1/aes_core/SB1/n2019 ), .Y(
        \U1/aes_core/SB1/n1814 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1293  ( .A(\U1/aes_core/SB1/n2017 ), .B(
        \U1/aes_core/SB1/n3346 ), .Y(\U1/aes_core/SB1/n2018 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1292  ( .A0(\U1/aes_core/SB1/n3331 ), 
        .A1(\U1/aes_core/SB1/n2018 ), .B0(\U1/aes_core/SB1/n3268 ), .Y(
        \U1/aes_core/SB1/n1813 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1291  ( .A0(\U1/aes_core/SB1/n2058 ), 
        .A1(\U1/aes_core/SB1/n3333 ), .B0(\U1/aes_core/SB1/n2055 ), .Y(
        \U1/aes_core/SB1/n1812 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1290  ( .A(\U1/aes_core/SB1/n2054 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n1851 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1289  ( .A(\U1/aes_core/SB1/n1814 ), .B(
        \U1/aes_core/SB1/n1813 ), .C(\U1/aes_core/SB1/n1812 ), .D(
        \U1/aes_core/SB1/n1851 ), .Y(\U1/aes_core/SB1/n1817 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1288  ( .A(\U1/aes_core/SB1/n3275 ), .B(
        \U1/aes_core/SB1/n2060 ), .Y(\U1/aes_core/SB1/n2059 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1287  ( .A(\U1/aes_core/SB1/n2053 ), .B(
        \U1/aes_core/SB1/n1976 ), .Y(\U1/aes_core/SB1/n1815 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1286  ( .A0(\U1/aes_core/SB1/n2059 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n1815 ), .B1(
        \U1/aes_core/SB1/n2010 ), .C0(\U1/aes_core/SB1/n3302 ), .C1(
        \U1/aes_core/SB1/n3278 ), .Y(\U1/aes_core/SB1/n1816 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1285  ( .A(\U1/aes_core/SB1/n3353 ), .B(
        \U1/aes_core/SB1/n3295 ), .C(\U1/aes_core/SB1/n2074 ), .D(
        \U1/aes_core/SB1/n1818 ), .E(\U1/aes_core/SB1/n1817 ), .F(
        \U1/aes_core/SB1/n1816 ), .Y(\U1/aes_core/sb1 [10]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1284  ( .A(\U1/aes_core/SB1/n3347 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n2034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1283  ( .A(\U1/aes_core/SB1/n3330 ), .B(
        \U1/aes_core/SB1/n1952 ), .Y(\U1/aes_core/SB1/n2036 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1282  ( .AN(\U1/aes_core/SB1/n1821 ), 
        .B(\U1/aes_core/SB1/n1820 ), .C(\U1/aes_core/SB1/n1819 ), .D(
        \U1/aes_core/SB1/n2036 ), .Y(\U1/aes_core/SB1/n1826 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1281  ( .A(\U1/aes_core/SB1/n3324 ), .B(
        \U1/aes_core/SB1/n2055 ), .Y(\U1/aes_core/SB1/n1983 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1280  ( .A0(\U1/aes_core/SB1/n3269 ), 
        .A1(\U1/aes_core/SB1/n3268 ), .B0(\U1/aes_core/SB1/n3323 ), .Y(
        \U1/aes_core/SB1/n1822 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1279  ( .A(\U1/aes_core/SB1/n3340 ), .B(
        \U1/aes_core/SB1/n1952 ), .Y(\U1/aes_core/SB1/n2061 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U1278  ( .A0(\U1/aes_core/SB1/n1983 ), 
        .A1(\U1/aes_core/SB1/n3296 ), .B0(\U1/aes_core/SB1/n1822 ), .C0(
        \U1/aes_core/SB1/n2061 ), .Y(\U1/aes_core/SB1/n1825 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1277  ( .A0(\U1/aes_core/SB1/n2020 ), 
        .A1(\U1/aes_core/SB1/n2070 ), .B0(\U1/aes_core/SB1/n1823 ), .B1(
        \U1/aes_core/SB1/n3308 ), .C0(\U1/aes_core/SB1/n3281 ), .C1(
        \U1/aes_core/SB1/n2065 ), .Y(\U1/aes_core/SB1/n1824 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1276  ( .A(\U1/aes_core/SB1/n1828 ), .B(
        \U1/aes_core/SB1/n2034 ), .C(\U1/aes_core/SB1/n1827 ), .D(
        \U1/aes_core/SB1/n1826 ), .E(\U1/aes_core/SB1/n1825 ), .F(
        \U1/aes_core/SB1/n1824 ), .Y(\U1/aes_core/SB1/n1962 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1275  ( .A(\U1/aes_core/SB1/n3323 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n2040 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1274  ( .AN(\U1/aes_core/SB1/n1831 ), 
        .B(\U1/aes_core/SB1/n1830 ), .C(\U1/aes_core/SB1/n1829 ), .D(
        \U1/aes_core/SB1/n2040 ), .Y(\U1/aes_core/SB1/n1838 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U1273  ( .A0(\U1/aes_core/SB1/n3331 ), 
        .A1(\U1/aes_core/SB1/n3327 ), .B0(\U1/aes_core/SB1/n3332 ), .B1(
        \U1/aes_core/SB1/n3334 ), .C0(\U1/aes_core/SB1/n3274 ), .C1(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n1837 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1272  ( .A0(\U1/aes_core/SB1/n3301 ), 
        .A1(\U1/aes_core/SB1/n3280 ), .B0(\U1/aes_core/SB1/n2021 ), .B1(
        \U1/aes_core/SB1/n2020 ), .Y(\U1/aes_core/SB1/n1832 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1271  ( .A0(\U1/aes_core/SB1/n1952 ), 
        .A1(\U1/aes_core/SB1/n3323 ), .B0(\U1/aes_core/SB1/n3276 ), .B1(
        \U1/aes_core/SB1/n3299 ), .C0(\U1/aes_core/SB1/n1832 ), .Y(
        \U1/aes_core/SB1/n1836 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1270  ( .A(\U1/aes_core/SB1/n3308 ), .B(
        \U1/aes_core/SB1/n3343 ), .Y(\U1/aes_core/SB1/n3270 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1269  ( .A(\U1/aes_core/SB1/n3344 ), .B(
        \U1/aes_core/SB1/n3347 ), .Y(\U1/aes_core/SB1/n1834 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1268  ( .A0(\U1/aes_core/SB1/n3340 ), 
        .A1(\U1/aes_core/SB1/n3270 ), .B0(\U1/aes_core/SB1/n2058 ), .B1(
        \U1/aes_core/SB1/n1834 ), .C0(\U1/aes_core/SB1/n1833 ), .Y(
        \U1/aes_core/SB1/n1835 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1267  ( .AN(\U1/aes_core/SB1/n1838 ), 
        .B(\U1/aes_core/SB1/n1837 ), .C(\U1/aes_core/SB1/n1836 ), .D(
        \U1/aes_core/SB1/n1835 ), .Y(\U1/aes_core/SB1/n1988 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1266  ( .A(\U1/aes_core/SB1/n1995 ), .B(
        \U1/aes_core/SB1/n3302 ), .Y(\U1/aes_core/SB1/n2024 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1265  ( .A0(\U1/aes_core/SB1/n3303 ), 
        .A1(\U1/aes_core/SB1/n3302 ), .B0(\U1/aes_core/SB1/n1839 ), .Y(
        \U1/aes_core/SB1/n1849 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1264  ( .A0(\U1/aes_core/SB1/n2058 ), 
        .A1(\U1/aes_core/SB1/n3332 ), .B0(\U1/aes_core/SB1/n3275 ), .B1(
        \U1/aes_core/SB1/n3307 ), .Y(\U1/aes_core/SB1/n1840 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1263  ( .A0(\U1/aes_core/SB1/n3344 ), 
        .A1(\U1/aes_core/SB1/n2039 ), .B0(\U1/aes_core/SB1/n2057 ), .B1(
        \U1/aes_core/SB1/n3343 ), .C0(\U1/aes_core/SB1/n1840 ), .Y(
        \U1/aes_core/SB1/n1848 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1262  ( .A(\U1/aes_core/SB1/n1912 ), .B(
        \U1/aes_core/SB1/n3308 ), .Y(\U1/aes_core/SB1/n3292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1261  ( .A(\U1/aes_core/SB1/n3305 ), .B(
        \U1/aes_core/SB1/n3323 ), .Y(\U1/aes_core/SB1/n2037 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1260  ( .AN(\U1/aes_core/SB1/n3292 ), 
        .B(\U1/aes_core/SB1/n1842 ), .C(\U1/aes_core/SB1/n1841 ), .D(
        \U1/aes_core/SB1/n2037 ), .Y(\U1/aes_core/SB1/n1847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1259  ( .A(\U1/aes_core/SB1/n3280 ), .B(
        \U1/aes_core/SB1/n3297 ), .Y(\U1/aes_core/SB1/n2015 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1258  ( .AN(\U1/aes_core/SB1/n2015 ), 
        .B(\U1/aes_core/SB1/n1845 ), .C(\U1/aes_core/SB1/n1844 ), .D(
        \U1/aes_core/SB1/n1843 ), .Y(\U1/aes_core/SB1/n1846 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1257  ( .A(\U1/aes_core/SB1/n2024 ), .B(
        \U1/aes_core/SB1/n1850 ), .C(\U1/aes_core/SB1/n1849 ), .D(
        \U1/aes_core/SB1/n1848 ), .E(\U1/aes_core/SB1/n1847 ), .F(
        \U1/aes_core/SB1/n1846 ), .Y(\U1/aes_core/SB1/n1924 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1256  ( .A(\U1/aes_core/SB1/n2017 ), .B(
        \U1/aes_core/SB1/n3300 ), .Y(\U1/aes_core/SB1/n2064 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1255  ( .A0(\U1/aes_core/SB1/n2017 ), 
        .A1(\U1/aes_core/SB1/n3280 ), .B0(\U1/aes_core/SB1/n1851 ), .Y(
        \U1/aes_core/SB1/n1861 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1254  ( .A(\U1/aes_core/SB1/n3343 ), .B(
        \U1/aes_core/SB1/n1912 ), .Y(\U1/aes_core/SB1/n2023 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1253  ( .A(\U1/aes_core/SB1/n1949 ), .B(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n3312 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1252  ( .AN(\U1/aes_core/SB1/n2023 ), 
        .B(\U1/aes_core/SB1/n1853 ), .C(\U1/aes_core/SB1/n1852 ), .D(
        \U1/aes_core/SB1/n3312 ), .Y(\U1/aes_core/SB1/n1860 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1251  ( .A(\U1/aes_core/SB1/n3274 ), .B(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n2045 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1250  ( .A(\U1/aes_core/SB1/n3339 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n3267 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1249  ( .A(\U1/aes_core/SB1/n2019 ), .B(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n3335 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1248  ( .A(\U1/aes_core/SB1/n1854 ), .B(
        \U1/aes_core/SB1/n2045 ), .C(\U1/aes_core/SB1/n3267 ), .D(
        \U1/aes_core/SB1/n3335 ), .Y(\U1/aes_core/SB1/n1859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1247  ( .A(\U1/aes_core/SB1/n3322 ), .B(
        \U1/aes_core/SB1/n3333 ), .Y(\U1/aes_core/SB1/n2005 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1246  ( .A(\U1/aes_core/SB1/n1857 ), .B(
        \U1/aes_core/SB1/n1856 ), .C(\U1/aes_core/SB1/n2005 ), .D(
        \U1/aes_core/SB1/n1855 ), .Y(\U1/aes_core/SB1/n1858 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1245  ( .A(\U1/aes_core/SB1/n2064 ), .B(
        \U1/aes_core/SB1/n1862 ), .C(\U1/aes_core/SB1/n1861 ), .D(
        \U1/aes_core/SB1/n1860 ), .E(\U1/aes_core/SB1/n1859 ), .F(
        \U1/aes_core/SB1/n1858 ), .Y(\U1/aes_core/SB1/n1940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1244  ( .A(\U1/aes_core/SB1/n3302 ), .B(
        \U1/aes_core/SB1/n2021 ), .Y(\U1/aes_core/SB1/n2016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1243  ( .A(\U1/aes_core/SB1/n3324 ), .B(
        \U1/aes_core/SB1/n3331 ), .Y(\U1/aes_core/SB1/n2041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1242  ( .A(\U1/aes_core/SB1/n3334 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n3265 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1241  ( .A(\U1/aes_core/SB1/n1864 ), .B(
        \U1/aes_core/SB1/n1863 ), .C(\U1/aes_core/SB1/n2041 ), .D(
        \U1/aes_core/SB1/n3265 ), .Y(\U1/aes_core/SB1/n1871 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1240  ( .A(\U1/aes_core/SB1/n1952 ), .B(
        \U1/aes_core/SB1/n3276 ), .Y(\U1/aes_core/SB1/n2027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1239  ( .A(\U1/aes_core/SB1/n3333 ), .B(
        \U1/aes_core/SB1/n1952 ), .Y(\U1/aes_core/SB1/n3311 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1238  ( .A(\U1/aes_core/SB1/n1866 ), .B(
        \U1/aes_core/SB1/n2027 ), .C(\U1/aes_core/SB1/n1865 ), .D(
        \U1/aes_core/SB1/n3311 ), .Y(\U1/aes_core/SB1/n1870 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U1237  ( .A(\U1/aes_core/SB1/n2055 ), .B(
        \U1/aes_core/SB1/n3329 ), .C(\U1/aes_core/SB1/n2053 ), .Y(
        \U1/aes_core/SB1/n1868 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1236  ( .A0(\U1/aes_core/SB1/n1868 ), 
        .A1(\U1/aes_core/SB1/n2010 ), .B0(\U1/aes_core/SB1/n2020 ), .B1(
        \U1/aes_core/SB1/n3347 ), .C0(\U1/aes_core/SB1/n1867 ), .Y(
        \U1/aes_core/SB1/n1869 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1235  ( .A(\U1/aes_core/SB1/n2016 ), .B(
        \U1/aes_core/SB1/n1873 ), .C(\U1/aes_core/SB1/n1872 ), .D(
        \U1/aes_core/SB1/n1871 ), .E(\U1/aes_core/SB1/n1870 ), .F(
        \U1/aes_core/SB1/n1869 ), .Y(\U1/aes_core/SB1/n1973 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1234  ( .A(\U1/aes_core/SB1/n3300 ), .B(
        \U1/aes_core/SB1/n1888 ), .Y(\U1/aes_core/SB1/n2028 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1233  ( .A0(\U1/aes_core/SB1/n2020 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n1874 ), .Y(
        \U1/aes_core/SB1/n1885 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1232  ( .A0(\U1/aes_core/SB1/n1976 ), 
        .A1(\U1/aes_core/SB1/n2019 ), .B0(\U1/aes_core/SB1/n3322 ), .B1(
        \U1/aes_core/SB1/n3334 ), .Y(\U1/aes_core/SB1/n1875 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1231  ( .A0(\U1/aes_core/SB1/n3308 ), 
        .A1(\U1/aes_core/SB1/n3346 ), .B0(\U1/aes_core/SB1/n3303 ), .B1(
        \U1/aes_core/SB1/n3279 ), .C0(\U1/aes_core/SB1/n1875 ), .Y(
        \U1/aes_core/SB1/n1884 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1230  ( .A(\U1/aes_core/SB1/n3303 ), .B(
        \U1/aes_core/SB1/n2020 ), .Y(\U1/aes_core/SB1/n3291 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1229  ( .A(\U1/aes_core/SB1/n3291 ), .Y(
        \U1/aes_core/SB1/n1877 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1228  ( .A(\U1/aes_core/SB1/n3332 ), .B(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n2047 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1227  ( .AN(\U1/aes_core/SB1/n1878 ), 
        .B(\U1/aes_core/SB1/n1877 ), .C(\U1/aes_core/SB1/n1876 ), .D(
        \U1/aes_core/SB1/n2047 ), .Y(\U1/aes_core/SB1/n1883 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1226  ( .A(\U1/aes_core/SB1/n2058 ), .B(
        \U1/aes_core/SB1/n3307 ), .Y(\U1/aes_core/SB1/n2003 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1225  ( .AN(\U1/aes_core/SB1/n1881 ), 
        .B(\U1/aes_core/SB1/n1880 ), .C(\U1/aes_core/SB1/n1879 ), .D(
        \U1/aes_core/SB1/n2003 ), .Y(\U1/aes_core/SB1/n1882 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1224  ( .A(\U1/aes_core/SB1/n2028 ), .B(
        \U1/aes_core/SB1/n1886 ), .C(\U1/aes_core/SB1/n1885 ), .D(
        \U1/aes_core/SB1/n1884 ), .E(\U1/aes_core/SB1/n1883 ), .F(
        \U1/aes_core/SB1/n1882 ), .Y(\U1/aes_core/SB1/n1947 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1223  ( .A0(\U1/aes_core/SB1/n2053 ), 
        .A1(\U1/aes_core/SB1/n2018 ), .B0(\U1/aes_core/SB1/n1976 ), .B1(
        \U1/aes_core/SB1/n2060 ), .Y(\U1/aes_core/SB1/n1887 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1222  ( .A0(\U1/aes_core/SB1/n3281 ), 
        .A1(\U1/aes_core/SB1/n3280 ), .B0(\U1/aes_core/SB1/n1888 ), .B1(
        \U1/aes_core/SB1/n3343 ), .C0(\U1/aes_core/SB1/n1887 ), .Y(
        \U1/aes_core/SB1/n1898 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1221  ( .A(\U1/aes_core/SB1/n3329 ), .B(
        \U1/aes_core/SB1/n3325 ), .Y(\U1/aes_core/SB1/n2044 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1220  ( .AN(\U1/aes_core/SB1/n1891 ), 
        .B(\U1/aes_core/SB1/n1890 ), .C(\U1/aes_core/SB1/n1889 ), .D(
        \U1/aes_core/SB1/n2044 ), .Y(\U1/aes_core/SB1/n1897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1219  ( .A0(\U1/aes_core/SB1/n3282 ), 
        .A1(\U1/aes_core/SB1/n3340 ), .B0(\U1/aes_core/SB1/n3322 ), .Y(
        \U1/aes_core/SB1/n1894 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1218  ( .A(\U1/aes_core/SB1/n3344 ), .B(
        \U1/aes_core/SB1/n1995 ), .Y(\U1/aes_core/SB1/n1892 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1217  ( .A0(\U1/aes_core/SB1/n3333 ), 
        .A1(\U1/aes_core/SB1/n1892 ), .B0(\U1/aes_core/SB1/n3329 ), .B1(
        \U1/aes_core/SB1/n1948 ), .Y(\U1/aes_core/SB1/n1893 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1216  ( .AN(\U1/aes_core/SB1/n1895 ), 
        .B(\U1/aes_core/SB1/n1894 ), .C(\U1/aes_core/SB1/n1893 ), .Y(
        \U1/aes_core/SB1/n1896 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1215  ( .A(\U1/aes_core/SB1/n1940 ), .B(
        \U1/aes_core/SB1/n1973 ), .C(\U1/aes_core/SB1/n1947 ), .D(
        \U1/aes_core/SB1/n1898 ), .E(\U1/aes_core/SB1/n1897 ), .F(
        \U1/aes_core/SB1/n1896 ), .Y(\U1/aes_core/SB1/n1999 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1214  ( .A(\U1/aes_core/SB1/n1962 ), .B(
        \U1/aes_core/SB1/n1988 ), .C(\U1/aes_core/SB1/n1924 ), .D(
        \U1/aes_core/SB1/n1999 ), .Y(\U1/aes_core/SB1/n1908 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1213  ( .A(\U1/aes_core/SB1/n3333 ), .B(
        \U1/aes_core/SB1/n2068 ), .Y(\U1/aes_core/SB1/n2009 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1212  ( .A(\U1/aes_core/SB1/n3323 ), .B(
        \U1/aes_core/SB1/n2060 ), .Y(\U1/aes_core/SB1/n2002 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1211  ( .A(\U1/aes_core/SB1/n3297 ), .B(
        \U1/aes_core/SB1/n3302 ), .Y(\U1/aes_core/SB1/n3306 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1210  ( .A0(\U1/aes_core/SB1/n1952 ), 
        .A1(\U1/aes_core/SB1/n3275 ), .B0(\U1/aes_core/SB1/n3306 ), .B1(
        \U1/aes_core/SB1/n3305 ), .Y(\U1/aes_core/SB1/n1899 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1209  ( .A0(\U1/aes_core/SB1/n2021 ), 
        .A1(\U1/aes_core/SB1/n2009 ), .B0(\U1/aes_core/SB1/n3278 ), .B1(
        \U1/aes_core/SB1/n2002 ), .C0(\U1/aes_core/SB1/n1899 ), .Y(
        \U1/aes_core/SB1/n1900 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1208  ( .A(\U1/aes_core/SB1/n1900 ), .Y(
        \U1/aes_core/SB1/n1907 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1207  ( .A0(\U1/aes_core/SB1/n3301 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n2020 ), .B1(
        \U1/aes_core/SB1/n1995 ), .Y(\U1/aes_core/SB1/n1901 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1206  ( .A0(\U1/aes_core/SB1/n2054 ), 
        .A1(\U1/aes_core/SB1/n3268 ), .B0(\U1/aes_core/SB1/n3327 ), .B1(
        \U1/aes_core/SB1/n3282 ), .C0(\U1/aes_core/SB1/n1901 ), .Y(
        \U1/aes_core/SB1/n1906 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1205  ( .A0(\U1/aes_core/SB1/n2068 ), 
        .A1(\U1/aes_core/SB1/n3323 ), .B0(\U1/aes_core/SB1/n2055 ), .Y(
        \U1/aes_core/SB1/n1904 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1204  ( .A(\U1/aes_core/SB1/n3340 ), .B(
        \U1/aes_core/SB1/n3305 ), .Y(\U1/aes_core/SB1/n2026 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB1/U1203  ( .A(\U1/aes_core/SB1/n1904 ), .B(
        \U1/aes_core/SB1/n2026 ), .C(\U1/aes_core/SB1/n1903 ), .D(
        \U1/aes_core/SB1/n1902 ), .Y(\U1/aes_core/SB1/n1905 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1202  ( .AN(\U1/aes_core/SB1/n1908 ), 
        .B(\U1/aes_core/SB1/n1907 ), .C(\U1/aes_core/SB1/n1906 ), .D(
        \U1/aes_core/SB1/n1905 ), .Y(\U1/aes_core/sb1 [11]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1201  ( .A0(\U1/aes_core/SB1/n1920 ), 
        .A1(\U1/aes_core/SB1/n2008 ), .B0(\U1/aes_core/SB1/n3297 ), .Y(
        \U1/aes_core/SB1/n1917 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1200  ( .A(\U1/aes_core/SB1/n1949 ), .B(
        \U1/aes_core/SB1/n3325 ), .Y(\U1/aes_core/SB1/n2035 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U1199  ( .A(\U1/aes_core/SB1/n1910 ), .B(
        \U1/aes_core/SB1/n2035 ), .C(\U1/aes_core/SB1/n1909 ), .Y(
        \U1/aes_core/SB1/n1916 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1198  ( .A(\U1/aes_core/SB1/n2053 ), .B(
        \U1/aes_core/SB1/n3322 ), .Y(\U1/aes_core/SB1/n1913 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1197  ( .A(\U1/aes_core/SB1/n3305 ), .B(
        \U1/aes_core/SB1/n1952 ), .Y(\U1/aes_core/SB1/n1911 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1196  ( .A0(\U1/aes_core/SB1/n1913 ), 
        .A1(\U1/aes_core/SB1/n1912 ), .B0(\U1/aes_core/SB1/n1911 ), .B1(
        \U1/aes_core/SB1/n2057 ), .C0(\U1/aes_core/SB1/n2006 ), .C1(
        \U1/aes_core/SB1/n2008 ), .Y(\U1/aes_core/SB1/n1915 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1195  ( .A0(\U1/aes_core/SB1/n3303 ), 
        .A1(\U1/aes_core/SB1/n2017 ), .B0(\U1/aes_core/SB1/n3281 ), .B1(
        \U1/aes_core/SB1/n3343 ), .C0(\U1/aes_core/SB1/n3308 ), .C1(
        \U1/aes_core/SB1/n2010 ), .Y(\U1/aes_core/SB1/n1914 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1194  ( .A(\U1/aes_core/SB1/n1919 ), .B(
        \U1/aes_core/SB1/n1918 ), .C(\U1/aes_core/SB1/n1917 ), .D(
        \U1/aes_core/SB1/n1916 ), .E(\U1/aes_core/SB1/n1915 ), .F(
        \U1/aes_core/SB1/n1914 ), .Y(\U1/aes_core/SB1/n2000 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1193  ( .A0(\U1/aes_core/SB1/n1920 ), 
        .A1(\U1/aes_core/SB1/n3280 ), .B0(\U1/aes_core/SB1/n3346 ), .Y(
        \U1/aes_core/SB1/n1946 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB1/U1192  ( .A0(\U1/aes_core/SB1/n3296 ), 
        .A1(\U1/aes_core/SB1/n3279 ), .A2(\U1/aes_core/SB1/n2010 ), .B0(
        \U1/aes_core/SB1/n3309 ), .Y(\U1/aes_core/SB1/n1945 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1191  ( .A(\U1/aes_core/SB1/n3276 ), .B(
        \U1/aes_core/SB1/n3327 ), .Y(\U1/aes_core/SB1/n2042 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1190  ( .A(\U1/aes_core/SB1/n1923 ), .B(
        \U1/aes_core/SB1/n1922 ), .C(\U1/aes_core/SB1/n1921 ), .D(
        \U1/aes_core/SB1/n2042 ), .Y(\U1/aes_core/SB1/n1942 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1189  ( .A(\U1/aes_core/SB1/n1924 ), .Y(
        \U1/aes_core/SB1/n1939 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1188  ( .A(\U1/aes_core/SB1/n3309 ), .B(
        \U1/aes_core/SB1/n3302 ), .Y(\U1/aes_core/SB1/n2022 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1187  ( .A0(\U1/aes_core/SB1/n2002 ), 
        .A1(\U1/aes_core/SB1/n2065 ), .B0(\U1/aes_core/SB1/n1925 ), .Y(
        \U1/aes_core/SB1/n1934 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1186  ( .A0(\U1/aes_core/SB1/n3280 ), 
        .A1(\U1/aes_core/SB1/n3342 ), .B0(\U1/aes_core/SB1/n3297 ), .B1(
        \U1/aes_core/SB1/n1995 ), .C0(\U1/aes_core/SB1/n3281 ), .C1(
        \U1/aes_core/SB1/n3309 ), .Y(\U1/aes_core/SB1/n1933 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1185  ( .A(\U1/aes_core/SB1/n3307 ), .B(
        \U1/aes_core/SB1/n3323 ), .Y(\U1/aes_core/SB1/n2046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1184  ( .A(\U1/aes_core/SB1/n2068 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n3272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1183  ( .A(\U1/aes_core/SB1/n1927 ), .B(
        \U1/aes_core/SB1/n1926 ), .C(\U1/aes_core/SB1/n2046 ), .D(
        \U1/aes_core/SB1/n3272 ), .Y(\U1/aes_core/SB1/n1932 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1182  ( .A(\U1/aes_core/SB1/n3333 ), .B(
        \U1/aes_core/SB1/n3299 ), .Y(\U1/aes_core/SB1/n2004 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1181  ( .AN(\U1/aes_core/SB1/n1930 ), 
        .B(\U1/aes_core/SB1/n1929 ), .C(\U1/aes_core/SB1/n1928 ), .D(
        \U1/aes_core/SB1/n2004 ), .Y(\U1/aes_core/SB1/n1931 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1180  ( .A(\U1/aes_core/SB1/n2022 ), .B(
        \U1/aes_core/SB1/n1935 ), .C(\U1/aes_core/SB1/n1934 ), .D(
        \U1/aes_core/SB1/n1933 ), .E(\U1/aes_core/SB1/n1932 ), .F(
        \U1/aes_core/SB1/n1931 ), .Y(\U1/aes_core/SB1/n1936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1179  ( .A(\U1/aes_core/SB1/n1936 ), .Y(
        \U1/aes_core/SB1/n1989 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1178  ( .A0(\U1/aes_core/SB1/n3344 ), 
        .A1(\U1/aes_core/SB1/n2017 ), .B0(\U1/aes_core/SB1/n3281 ), .B1(
        \U1/aes_core/SB1/n3347 ), .Y(\U1/aes_core/SB1/n1937 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U1177  ( .A0(\U1/aes_core/SB1/n3324 ), 
        .A1(\U1/aes_core/SB1/n3323 ), .B0(\U1/aes_core/SB1/n3330 ), .B1(
        \U1/aes_core/SB1/n3299 ), .C0(\U1/aes_core/SB1/n1937 ), .Y(
        \U1/aes_core/SB1/n1938 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1176  ( .AN(\U1/aes_core/SB1/n1940 ), 
        .B(\U1/aes_core/SB1/n1939 ), .C(\U1/aes_core/SB1/n1989 ), .D(
        \U1/aes_core/SB1/n1938 ), .Y(\U1/aes_core/SB1/n1941 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1175  ( .A(\U1/aes_core/SB1/n1946 ), .B(
        \U1/aes_core/SB1/n1945 ), .C(\U1/aes_core/SB1/n1944 ), .D(
        \U1/aes_core/SB1/n1943 ), .E(\U1/aes_core/SB1/n1942 ), .F(
        \U1/aes_core/SB1/n1941 ), .Y(\U1/aes_core/SB1/n1987 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1174  ( .A(\U1/aes_core/SB1/n1947 ), .Y(
        \U1/aes_core/SB1/n1951 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1173  ( .A0(\U1/aes_core/SB1/n1949 ), 
        .A1(\U1/aes_core/SB1/n1948 ), .B0(\U1/aes_core/SB1/n1952 ), .B1(
        \U1/aes_core/SB1/n3339 ), .Y(\U1/aes_core/SB1/n1950 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U1172  ( .A0(\U1/aes_core/SB1/n2006 ), 
        .A1(\U1/aes_core/SB1/n3309 ), .B0(\U1/aes_core/SB1/n1951 ), .C0(
        \U1/aes_core/SB1/n1950 ), .Y(\U1/aes_core/SB1/n1961 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1171  ( .A0(\U1/aes_core/SB1/n3276 ), 
        .A1(\U1/aes_core/SB1/n3275 ), .B0(\U1/aes_core/SB1/n3332 ), .Y(
        \U1/aes_core/SB1/n1956 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1170  ( .A0(\U1/aes_core/SB1/n1952 ), 
        .A1(\U1/aes_core/SB1/n3268 ), .B0(\U1/aes_core/SB1/n2060 ), .Y(
        \U1/aes_core/SB1/n1955 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1169  ( .A(\U1/aes_core/SB1/n1956 ), .B(
        \U1/aes_core/SB1/n1955 ), .C(\U1/aes_core/SB1/n1954 ), .D(
        \U1/aes_core/SB1/n1953 ), .Y(\U1/aes_core/SB1/n1960 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1168  ( .A(\U1/aes_core/SB1/n3325 ), .B(
        \U1/aes_core/SB1/n3334 ), .Y(\U1/aes_core/SB1/n1958 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1167  ( .A(\U1/aes_core/SB1/n3331 ), .B(
        \U1/aes_core/SB1/n3333 ), .Y(\U1/aes_core/SB1/n1957 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1166  ( .A(\U1/aes_core/SB1/n1976 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n3310 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1165  ( .A0(\U1/aes_core/SB1/n1958 ), 
        .A1(\U1/aes_core/SB1/n2070 ), .B0(\U1/aes_core/SB1/n1957 ), .B1(
        \U1/aes_core/SB1/n2008 ), .C0(\U1/aes_core/SB1/n3310 ), .C1(
        \U1/aes_core/SB1/n2039 ), .Y(\U1/aes_core/SB1/n1959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1164  ( .A(\U1/aes_core/SB1/n2000 ), .B(
        \U1/aes_core/SB1/n1987 ), .C(\U1/aes_core/SB1/n1962 ), .D(
        \U1/aes_core/SB1/n1961 ), .E(\U1/aes_core/SB1/n1960 ), .F(
        \U1/aes_core/SB1/n1959 ), .Y(\U1/aes_core/sb1 [12]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1163  ( .A(\U1/aes_core/SB1/n3300 ), .B(
        \U1/aes_core/SB1/n3297 ), .Y(\U1/aes_core/SB1/n2025 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U1162  ( .A1N(\U1/aes_core/SB1/n3306 ), 
        .A0(\U1/aes_core/SB1/n3279 ), .B0(\U1/aes_core/SB1/n3344 ), .Y(
        \U1/aes_core/SB1/n1971 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1161  ( .A(\U1/aes_core/SB1/n2053 ), .B(
        \U1/aes_core/SB1/n3268 ), .Y(\U1/aes_core/SB1/n1963 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1160  ( .A0(\U1/aes_core/SB1/n2070 ), 
        .A1(\U1/aes_core/SB1/n3302 ), .B0(\U1/aes_core/SB1/n1963 ), .B1(
        \U1/aes_core/SB1/n3281 ), .C0(\U1/aes_core/SB1/n3297 ), .C1(
        \U1/aes_core/SB1/n3278 ), .Y(\U1/aes_core/SB1/n1970 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1159  ( .A(\U1/aes_core/SB1/n3327 ), .B(
        \U1/aes_core/SB1/n2019 ), .Y(\U1/aes_core/SB1/n2043 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1158  ( .A(\U1/aes_core/SB1/n3299 ), .B(
        \U1/aes_core/SB1/n3282 ), .Y(\U1/aes_core/SB1/n3266 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1157  ( .AN(\U1/aes_core/SB1/n1965 ), 
        .B(\U1/aes_core/SB1/n1964 ), .C(\U1/aes_core/SB1/n2043 ), .D(
        \U1/aes_core/SB1/n3266 ), .Y(\U1/aes_core/SB1/n1969 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1156  ( .A(\U1/aes_core/SB1/n3269 ), .B(
        \U1/aes_core/SB1/n3330 ), .Y(\U1/aes_core/SB1/n3313 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1155  ( .AN(\U1/aes_core/SB1/n1967 ), 
        .B(\U1/aes_core/SB1/n1966 ), .C(\U1/aes_core/SB1/n3313 ), .Y(
        \U1/aes_core/SB1/n1968 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1154  ( .A(\U1/aes_core/SB1/n2025 ), .B(
        \U1/aes_core/SB1/n1972 ), .C(\U1/aes_core/SB1/n1971 ), .D(
        \U1/aes_core/SB1/n1970 ), .E(\U1/aes_core/SB1/n1969 ), .F(
        \U1/aes_core/SB1/n1968 ), .Y(\U1/aes_core/SB1/n2001 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1153  ( .A(\U1/aes_core/SB1/n1973 ), .Y(
        \U1/aes_core/SB1/n1975 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1152  ( .A0(\U1/aes_core/SB1/n3322 ), 
        .A1(\U1/aes_core/SB1/n2058 ), .B0(\U1/aes_core/SB1/n2060 ), .B1(
        \U1/aes_core/SB1/n3327 ), .Y(\U1/aes_core/SB1/n1974 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U1151  ( .A0(\U1/aes_core/SB1/n3344 ), 
        .A1(\U1/aes_core/SB1/n3346 ), .B0(\U1/aes_core/SB1/n1975 ), .C0(
        \U1/aes_core/SB1/n1974 ), .Y(\U1/aes_core/SB1/n1986 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1150  ( .A0(\U1/aes_core/SB1/n3324 ), 
        .A1(\U1/aes_core/SB1/n3322 ), .B0(\U1/aes_core/SB1/n2019 ), .Y(
        \U1/aes_core/SB1/n1979 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1149  ( .A0(\U1/aes_core/SB1/n3325 ), 
        .A1(\U1/aes_core/SB1/n3339 ), .B0(\U1/aes_core/SB1/n1976 ), .Y(
        \U1/aes_core/SB1/n1978 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1148  ( .AN(\U1/aes_core/SB1/n1980 ), 
        .B(\U1/aes_core/SB1/n1979 ), .C(\U1/aes_core/SB1/n1978 ), .D(
        \U1/aes_core/SB1/n1977 ), .Y(\U1/aes_core/SB1/n1985 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1147  ( .A0(\U1/aes_core/SB1/n3332 ), 
        .A1(\U1/aes_core/SB1/n3329 ), .B0(\U1/aes_core/SB1/n3333 ), .Y(
        \U1/aes_core/SB1/n1982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1146  ( .A(\U1/aes_core/SB1/n2017 ), .B(
        \U1/aes_core/SB1/n3302 ), .Y(\U1/aes_core/SB1/n3341 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1145  ( .A0(\U1/aes_core/SB1/n3307 ), 
        .A1(\U1/aes_core/SB1/n3341 ), .B0(\U1/aes_core/SB1/n2054 ), .B1(
        \U1/aes_core/SB1/n3305 ), .Y(\U1/aes_core/SB1/n1981 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U1144  ( .A0(\U1/aes_core/SB1/n1983 ), 
        .A1(\U1/aes_core/SB1/n2039 ), .B0(\U1/aes_core/SB1/n1982 ), .C0(
        \U1/aes_core/SB1/n1981 ), .Y(\U1/aes_core/SB1/n1984 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1143  ( .A(\U1/aes_core/SB1/n2001 ), .B(
        \U1/aes_core/SB1/n1988 ), .C(\U1/aes_core/SB1/n1987 ), .D(
        \U1/aes_core/SB1/n1986 ), .E(\U1/aes_core/SB1/n1985 ), .F(
        \U1/aes_core/SB1/n1984 ), .Y(\U1/aes_core/sb1 [13]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1142  ( .A0(\U1/aes_core/SB1/n3343 ), 
        .A1(\U1/aes_core/SB1/n3296 ), .B0(\U1/aes_core/SB1/n3301 ), .B1(
        \U1/aes_core/SB1/n2070 ), .C0(\U1/aes_core/SB1/n1989 ), .Y(
        \U1/aes_core/SB1/n1998 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1141  ( .A0(\U1/aes_core/SB1/n3275 ), 
        .A1(\U1/aes_core/SB1/n2068 ), .B0(\U1/aes_core/SB1/n3322 ), .Y(
        \U1/aes_core/SB1/n1993 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1140  ( .A0(\U1/aes_core/SB1/n2055 ), 
        .A1(\U1/aes_core/SB1/n3299 ), .B0(\U1/aes_core/SB1/n2060 ), .Y(
        \U1/aes_core/SB1/n1992 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1139  ( .A(\U1/aes_core/SB1/n2010 ), .B(
        \U1/aes_core/SB1/n3346 ), .Y(\U1/aes_core/SB1/n3328 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1138  ( .A0(\U1/aes_core/SB1/n3305 ), 
        .A1(\U1/aes_core/SB1/n3268 ), .B0(\U1/aes_core/SB1/n3328 ), .Y(
        \U1/aes_core/SB1/n1991 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1137  ( .A(\U1/aes_core/SB1/n1993 ), .B(
        \U1/aes_core/SB1/n1992 ), .C(\U1/aes_core/SB1/n1991 ), .D(
        \U1/aes_core/SB1/n1990 ), .Y(\U1/aes_core/SB1/n1997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1136  ( .A(\U1/aes_core/SB1/n3343 ), .B(
        \U1/aes_core/SB1/n3344 ), .Y(\U1/aes_core/SB1/n2066 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1135  ( .A(\U1/aes_core/SB1/n3332 ), .B(
        \U1/aes_core/SB1/n2066 ), .Y(\U1/aes_core/SB1/n1994 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1134  ( .A0(\U1/aes_core/SB1/n2057 ), 
        .A1(\U1/aes_core/SB1/n1995 ), .B0(\U1/aes_core/SB1/n1994 ), .B1(
        \U1/aes_core/SB1/n2010 ), .C0(\U1/aes_core/SB1/n2008 ), .C1(
        \U1/aes_core/SB1/n2039 ), .Y(\U1/aes_core/SB1/n1996 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1133  ( .A(\U1/aes_core/SB1/n2001 ), .B(
        \U1/aes_core/SB1/n2000 ), .C(\U1/aes_core/SB1/n1999 ), .D(
        \U1/aes_core/SB1/n1998 ), .E(\U1/aes_core/SB1/n1997 ), .F(
        \U1/aes_core/SB1/n1996 ), .Y(\U1/aes_core/sb1 [14]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1132  ( .A0(\U1/aes_core/SB1/n2002 ), 
        .A1(\U1/aes_core/SB1/n3302 ), .B0(\U1/aes_core/SB1/n2070 ), .Y(
        \U1/aes_core/SB1/n2014 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U1131  ( .A(\U1/aes_core/SB1/n2005 ), .B(
        \U1/aes_core/SB1/n2004 ), .C(\U1/aes_core/SB1/n2003 ), .Y(
        \U1/aes_core/SB1/n2013 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U1130  ( .A(\U1/aes_core/SB1/n2054 ), .B(
        \U1/aes_core/SB1/n2058 ), .C(\U1/aes_core/SB1/n3282 ), .Y(
        \U1/aes_core/SB1/n2007 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1129  ( .A0(\U1/aes_core/SB1/n2009 ), 
        .A1(\U1/aes_core/SB1/n2008 ), .B0(\U1/aes_core/SB1/n2007 ), .B1(
        \U1/aes_core/SB1/n2065 ), .C0(\U1/aes_core/SB1/n2006 ), .C1(
        \U1/aes_core/SB1/n3280 ), .Y(\U1/aes_core/SB1/n2012 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U1128  ( .A0(\U1/aes_core/SB1/n3343 ), 
        .A1(\U1/aes_core/SB1/n2039 ), .B0(\U1/aes_core/SB1/n3344 ), .B1(
        \U1/aes_core/SB1/n2010 ), .Y(\U1/aes_core/SB1/n2011 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1127  ( .A(\U1/aes_core/SB1/n2016 ), .B(
        \U1/aes_core/SB1/n2015 ), .C(\U1/aes_core/SB1/n2014 ), .D(
        \U1/aes_core/SB1/n2013 ), .E(\U1/aes_core/SB1/n2012 ), .F(
        \U1/aes_core/SB1/n2011 ), .Y(\U1/aes_core/SB1/n3352 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U1126  ( .A0(\U1/aes_core/SB1/n3278 ), 
        .A1(\U1/aes_core/SB1/n3347 ), .B0(\U1/aes_core/SB1/n2017 ), .Y(
        \U1/aes_core/SB1/n2033 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB1/U1125  ( .A0(\U1/aes_core/SB1/n2019 ), 
        .A1(\U1/aes_core/SB1/n3269 ), .B0(\U1/aes_core/SB1/n2018 ), .B1(
        \U1/aes_core/SB1/n3329 ), .Y(\U1/aes_core/SB1/n2032 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1124  ( .A0(\U1/aes_core/SB1/n3281 ), 
        .A1(\U1/aes_core/SB1/n3344 ), .B0(\U1/aes_core/SB1/n2021 ), .B1(
        \U1/aes_core/SB1/n2020 ), .C0(\U1/aes_core/SB1/n2039 ), .C1(
        \U1/aes_core/SB1/n2065 ), .Y(\U1/aes_core/SB1/n2031 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1123  ( .A(\U1/aes_core/SB1/n2025 ), .B(
        \U1/aes_core/SB1/n2024 ), .C(\U1/aes_core/SB1/n2023 ), .D(
        \U1/aes_core/SB1/n2022 ), .Y(\U1/aes_core/SB1/n2030 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1122  ( .AN(\U1/aes_core/SB1/n2028 ), 
        .B(\U1/aes_core/SB1/n2027 ), .C(\U1/aes_core/SB1/n2026 ), .Y(
        \U1/aes_core/SB1/n2029 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1121  ( .A(\U1/aes_core/SB1/n2034 ), .B(
        \U1/aes_core/SB1/n2033 ), .C(\U1/aes_core/SB1/n2032 ), .D(
        \U1/aes_core/SB1/n2031 ), .E(\U1/aes_core/SB1/n2030 ), .F(
        \U1/aes_core/SB1/n2029 ), .Y(\U1/aes_core/SB1/n3294 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1120  ( .A0(\U1/aes_core/SB1/n3307 ), 
        .A1(\U1/aes_core/SB1/n3327 ), .B0(\U1/aes_core/SB1/n2054 ), .Y(
        \U1/aes_core/SB1/n2038 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1119  ( .A(\U1/aes_core/SB1/n2038 ), .B(
        \U1/aes_core/SB1/n2037 ), .C(\U1/aes_core/SB1/n2036 ), .D(
        \U1/aes_core/SB1/n2035 ), .Y(\U1/aes_core/SB1/n2051 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1118  ( .A0(\U1/aes_core/SB1/n3301 ), 
        .A1(\U1/aes_core/SB1/n2070 ), .B0(\U1/aes_core/SB1/n3279 ), .B1(
        \U1/aes_core/SB1/n3280 ), .C0(\U1/aes_core/SB1/n3309 ), .C1(
        \U1/aes_core/SB1/n2039 ), .Y(\U1/aes_core/SB1/n2050 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1117  ( .A(\U1/aes_core/SB1/n2043 ), .B(
        \U1/aes_core/SB1/n2042 ), .C(\U1/aes_core/SB1/n2041 ), .D(
        \U1/aes_core/SB1/n2040 ), .Y(\U1/aes_core/SB1/n2049 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U1116  ( .A(\U1/aes_core/SB1/n2047 ), .B(
        \U1/aes_core/SB1/n2046 ), .C(\U1/aes_core/SB1/n2045 ), .D(
        \U1/aes_core/SB1/n2044 ), .Y(\U1/aes_core/SB1/n2048 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1115  ( .A(\U1/aes_core/SB1/n2051 ), .B(
        \U1/aes_core/SB1/n2050 ), .C(\U1/aes_core/SB1/n2049 ), .D(
        \U1/aes_core/SB1/n2048 ), .Y(\U1/aes_core/SB1/n2052 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1114  ( .A(\U1/aes_core/SB1/n2052 ), .Y(
        \U1/aes_core/SB1/n3285 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1113  ( .A0(\U1/aes_core/SB1/n2055 ), 
        .A1(\U1/aes_core/SB1/n3330 ), .B0(\U1/aes_core/SB1/n2054 ), .B1(
        \U1/aes_core/SB1/n2053 ), .Y(\U1/aes_core/SB1/n2056 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U1112  ( .A0(\U1/aes_core/SB1/n2057 ), 
        .A1(\U1/aes_core/SB1/n3309 ), .B0(\U1/aes_core/SB1/n3285 ), .C0(
        \U1/aes_core/SB1/n2056 ), .Y(\U1/aes_core/SB1/n2073 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U1111  ( .A1N(\U1/aes_core/SB1/n2059 ), 
        .A0(\U1/aes_core/SB1/n2058 ), .B0(\U1/aes_core/SB1/n3332 ), .Y(
        \U1/aes_core/SB1/n2063 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1110  ( .A0(\U1/aes_core/SB1/n3327 ), 
        .A1(\U1/aes_core/SB1/n3322 ), .B0(\U1/aes_core/SB1/n2060 ), .Y(
        \U1/aes_core/SB1/n2062 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1109  ( .AN(\U1/aes_core/SB1/n2064 ), 
        .B(\U1/aes_core/SB1/n2063 ), .C(\U1/aes_core/SB1/n2062 ), .D(
        \U1/aes_core/SB1/n2061 ), .Y(\U1/aes_core/SB1/n2072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1108  ( .A(\U1/aes_core/SB1/n2065 ), .B(
        \U1/aes_core/SB1/n3343 ), .Y(\U1/aes_core/SB1/n2067 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1107  ( .A0(\U1/aes_core/SB1/n2068 ), 
        .A1(\U1/aes_core/SB1/n2067 ), .B0(\U1/aes_core/SB1/n3282 ), .B1(
        \U1/aes_core/SB1/n2066 ), .Y(\U1/aes_core/SB1/n2069 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1106  ( .A0(\U1/aes_core/SB1/n3281 ), 
        .A1(\U1/aes_core/SB1/n3347 ), .B0(\U1/aes_core/SB1/n2070 ), .B1(
        \U1/aes_core/SB1/n3342 ), .C0(\U1/aes_core/SB1/n2069 ), .Y(
        \U1/aes_core/SB1/n2071 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U1105  ( .A(\U1/aes_core/SB1/n3352 ), .B(
        \U1/aes_core/SB1/n3294 ), .C(\U1/aes_core/SB1/n2074 ), .D(
        \U1/aes_core/SB1/n2073 ), .E(\U1/aes_core/SB1/n2072 ), .F(
        \U1/aes_core/SB1/n2071 ), .Y(\U1/aes_core/sb1 [15]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1104  ( .A(Dout[87]), .B(Dout[86]), .Y(
        \U1/aes_core/SB1/n2093 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1103  ( .A(Dout[85]), .B(Dout[84]), .Y(
        \U1/aes_core/SB1/n2084 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1102  ( .A(\U1/aes_core/SB1/n2093 ), .B(
        \U1/aes_core/SB1/n2084 ), .Y(\U1/aes_core/SB1/n2157 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1101  ( .A(Dout[81]), .Y(
        \U1/aes_core/SB1/n2078 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1100  ( .A(Dout[80]), .Y(
        \U1/aes_core/SB1/n2075 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1099  ( .A(\U1/aes_core/SB1/n2078 ), .B(
        \U1/aes_core/SB1/n2075 ), .Y(\U1/aes_core/SB1/n2085 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1098  ( .A(Dout[83]), .B(Dout[82]), .Y(
        \U1/aes_core/SB1/n2105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1097  ( .A(\U1/aes_core/SB1/n2085 ), .B(
        \U1/aes_core/SB1/n2105 ), .Y(\U1/aes_core/SB1/n2464 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1096  ( .A(\U1/aes_core/SB1/n2157 ), .B(
        \U1/aes_core/SB1/n2464 ), .Y(\U1/aes_core/SB1/n2246 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U1095  ( .A(Dout[82]), .B(Dout[83]), .Y(
        \U1/aes_core/SB1/n2088 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1094  ( .A(\U1/aes_core/SB1/n2088 ), .B(
        \U1/aes_core/SB1/n2085 ), .Y(\U1/aes_core/SB1/n2402 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1093  ( .A(Dout[87]), .Y(
        \U1/aes_core/SB1/n2081 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1092  ( .A(\U1/aes_core/SB1/n2081 ), .B(
        Dout[86]), .Y(\U1/aes_core/SB1/n2111 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1091  ( .A(\U1/aes_core/SB1/n2111 ), .B(
        \U1/aes_core/SB1/n2084 ), .Y(\U1/aes_core/SB1/n2156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1090  ( .A(\U1/aes_core/SB1/n2402 ), .B(
        \U1/aes_core/SB1/n2156 ), .Y(\U1/aes_core/SB1/n2368 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1089  ( .A(Dout[83]), .Y(
        \U1/aes_core/SB1/n2076 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U1088  ( .A(Dout[82]), .B(
        \U1/aes_core/SB1/n2076 ), .Y(\U1/aes_core/SB1/n2086 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1087  ( .A(\U1/aes_core/SB1/n2085 ), .B(
        \U1/aes_core/SB1/n2086 ), .Y(\U1/aes_core/SB1/n2308 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1086  ( .A(\U1/aes_core/SB1/n2308 ), .Y(
        \U1/aes_core/SB1/n2498 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1085  ( .A(Dout[84]), .Y(
        \U1/aes_core/SB1/n2077 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1084  ( .A(\U1/aes_core/SB1/n2077 ), .B(
        Dout[85]), .Y(\U1/aes_core/SB1/n2092 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1083  ( .A(Dout[86]), .Y(
        \U1/aes_core/SB1/n2080 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1082  ( .A(\U1/aes_core/SB1/n2080 ), .B(
        Dout[87]), .Y(\U1/aes_core/SB1/n2102 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1081  ( .A(\U1/aes_core/SB1/n2092 ), .B(
        \U1/aes_core/SB1/n2102 ), .Y(\U1/aes_core/SB1/n2354 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1080  ( .A(\U1/aes_core/SB1/n2354 ), .Y(
        \U1/aes_core/SB1/n2452 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1079  ( .A(\U1/aes_core/SB1/n2498 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2286 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1078  ( .A(\U1/aes_core/SB1/n2157 ), .Y(
        \U1/aes_core/SB1/n2467 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1077  ( .A(Dout[81]), .B(Dout[80]), .Y(
        \U1/aes_core/SB1/n2089 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1076  ( .A(\U1/aes_core/SB1/n2089 ), .B(
        \U1/aes_core/SB1/n2105 ), .Y(\U1/aes_core/SB1/n2420 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1075  ( .A(\U1/aes_core/SB1/n2420 ), .Y(
        \U1/aes_core/SB1/n2508 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1074  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2508 ), .Y(\U1/aes_core/SB1/n2425 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1073  ( .A(\U1/aes_core/SB1/n2075 ), .B(
        Dout[81]), .Y(\U1/aes_core/SB1/n2104 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1072  ( .A(\U1/aes_core/SB1/n2086 ), .B(
        \U1/aes_core/SB1/n2104 ), .Y(\U1/aes_core/SB1/n2295 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1071  ( .A(\U1/aes_core/SB1/n2295 ), .Y(
        \U1/aes_core/SB1/n2409 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1070  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2264 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U1069  ( .A(\U1/aes_core/SB1/n2286 ), .B(
        \U1/aes_core/SB1/n2425 ), .C(\U1/aes_core/SB1/n2264 ), .Y(
        \U1/aes_core/SB1/n2124 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1068  ( .A(\U1/aes_core/SB1/n2084 ), .B(
        \U1/aes_core/SB1/n2102 ), .Y(\U1/aes_core/SB1/n2353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1067  ( .A(\U1/aes_core/SB1/n2076 ), .B(
        Dout[82]), .Y(\U1/aes_core/SB1/n2095 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1066  ( .A(\U1/aes_core/SB1/n2095 ), .B(
        \U1/aes_core/SB1/n2104 ), .Y(\U1/aes_core/SB1/n2351 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1065  ( .A(\U1/aes_core/SB1/n2353 ), .B(
        \U1/aes_core/SB1/n2351 ), .Y(\U1/aes_core/SB1/n2241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1064  ( .A(\U1/aes_core/SB1/n2156 ), .Y(
        \U1/aes_core/SB1/n2469 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1063  ( .A(Dout[85]), .Y(
        \U1/aes_core/SB1/n2079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1062  ( .A(\U1/aes_core/SB1/n2077 ), .B(
        \U1/aes_core/SB1/n2079 ), .Y(\U1/aes_core/SB1/n2103 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1061  ( .A(\U1/aes_core/SB1/n2093 ), .B(
        \U1/aes_core/SB1/n2103 ), .Y(\U1/aes_core/SB1/n2512 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1060  ( .A(\U1/aes_core/SB1/n2512 ), .Y(
        \U1/aes_core/SB1/n2443 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1059  ( .A(\U1/aes_core/SB1/n2078 ), .B(
        Dout[80]), .Y(\U1/aes_core/SB1/n2094 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1058  ( .A(\U1/aes_core/SB1/n2094 ), .B(
        \U1/aes_core/SB1/n2105 ), .Y(\U1/aes_core/SB1/n2477 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1057  ( .A(\U1/aes_core/SB1/n2477 ), .Y(
        \U1/aes_core/SB1/n2300 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1056  ( .A0(\U1/aes_core/SB1/n2469 ), 
        .A1(\U1/aes_core/SB1/n2443 ), .B0(\U1/aes_core/SB1/n2300 ), .Y(
        \U1/aes_core/SB1/n2083 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1055  ( .A(\U1/aes_core/SB1/n2089 ), .B(
        \U1/aes_core/SB1/n2086 ), .Y(\U1/aes_core/SB1/n2465 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1054  ( .A(\U1/aes_core/SB1/n2465 ), .Y(
        \U1/aes_core/SB1/n2451 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1053  ( .A(\U1/aes_core/SB1/n2079 ), .B(
        Dout[84]), .Y(\U1/aes_core/SB1/n2110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1052  ( .A(\U1/aes_core/SB1/n2102 ), .B(
        \U1/aes_core/SB1/n2110 ), .Y(\U1/aes_core/SB1/n2505 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1051  ( .A(\U1/aes_core/SB1/n2353 ), .B(
        \U1/aes_core/SB1/n2505 ), .Y(\U1/aes_core/SB1/n2219 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1050  ( .A(\U1/aes_core/SB1/n2081 ), .B(
        \U1/aes_core/SB1/n2080 ), .Y(\U1/aes_core/SB1/n2101 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1049  ( .A(\U1/aes_core/SB1/n2092 ), .B(
        \U1/aes_core/SB1/n2101 ), .Y(\U1/aes_core/SB1/n2480 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1048  ( .A(\U1/aes_core/SB1/n2480 ), .Y(
        \U1/aes_core/SB1/n2200 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1047  ( .A0(\U1/aes_core/SB1/n2451 ), 
        .A1(\U1/aes_core/SB1/n2219 ), .B0(\U1/aes_core/SB1/n2200 ), .B1(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2082 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U1046  ( .AN(\U1/aes_core/SB1/n2241 ), 
        .B(\U1/aes_core/SB1/n2083 ), .C(\U1/aes_core/SB1/n2082 ), .Y(
        \U1/aes_core/SB1/n2123 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1045  ( .A(\U1/aes_core/SB1/n2084 ), .B(
        \U1/aes_core/SB1/n2101 ), .Y(\U1/aes_core/SB1/n2370 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1044  ( .A(\U1/aes_core/SB1/n2088 ), .B(
        \U1/aes_core/SB1/n2089 ), .Y(\U1/aes_core/SB1/n2515 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1043  ( .A(\U1/aes_core/SB1/n2111 ), .B(
        \U1/aes_core/SB1/n2092 ), .Y(\U1/aes_core/SB1/n2421 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1042  ( .A(\U1/aes_core/SB1/n2088 ), .B(
        \U1/aes_core/SB1/n2094 ), .Y(\U1/aes_core/SB1/n2418 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1041  ( .A(\U1/aes_core/SB1/n2085 ), .B(
        \U1/aes_core/SB1/n2095 ), .Y(\U1/aes_core/SB1/n2423 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1040  ( .A(\U1/aes_core/SB1/n2423 ), .Y(
        \U1/aes_core/SB1/n2403 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1039  ( .A(\U1/aes_core/SB1/n2505 ), .Y(
        \U1/aes_core/SB1/n2214 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1038  ( .A(\U1/aes_core/SB1/n2086 ), .B(
        \U1/aes_core/SB1/n2094 ), .Y(\U1/aes_core/SB1/n2441 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1037  ( .A(\U1/aes_core/SB1/n2441 ), .Y(
        \U1/aes_core/SB1/n2466 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U1036  ( .A0(\U1/aes_core/SB1/n2403 ), 
        .A1(\U1/aes_core/SB1/n2467 ), .B0(\U1/aes_core/SB1/n2214 ), .B1(
        \U1/aes_core/SB1/n2466 ), .Y(\U1/aes_core/SB1/n2087 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U1035  ( .A0(\U1/aes_core/SB1/n2370 ), 
        .A1(\U1/aes_core/SB1/n2515 ), .B0(\U1/aes_core/SB1/n2421 ), .B1(
        \U1/aes_core/SB1/n2418 ), .C0(\U1/aes_core/SB1/n2087 ), .Y(
        \U1/aes_core/SB1/n2122 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1034  ( .A(\U1/aes_core/SB1/n2423 ), .B(
        \U1/aes_core/SB1/n2370 ), .Y(\U1/aes_core/SB1/n2207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1033  ( .A(\U1/aes_core/SB1/n2418 ), .B(
        \U1/aes_core/SB1/n2353 ), .Y(\U1/aes_core/SB1/n2217 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1032  ( .A(\U1/aes_core/SB1/n2217 ), .Y(
        \U1/aes_core/SB1/n2091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1031  ( .A(\U1/aes_core/SB1/n2088 ), .B(
        \U1/aes_core/SB1/n2104 ), .Y(\U1/aes_core/SB1/n2493 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1030  ( .A(\U1/aes_core/SB1/n2493 ), .Y(
        \U1/aes_core/SB1/n2442 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1029  ( .A(\U1/aes_core/SB1/n2089 ), .B(
        \U1/aes_core/SB1/n2095 ), .Y(\U1/aes_core/SB1/n2478 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1028  ( .A(\U1/aes_core/SB1/n2478 ), .Y(
        \U1/aes_core/SB1/n2489 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U1027  ( .A0(\U1/aes_core/SB1/n2442 ), 
        .A1(\U1/aes_core/SB1/n2489 ), .B0(\U1/aes_core/SB1/n2443 ), .Y(
        \U1/aes_core/SB1/n2090 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1026  ( .A(\U1/aes_core/SB1/n2093 ), .B(
        \U1/aes_core/SB1/n2110 ), .Y(\U1/aes_core/SB1/n2494 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1025  ( .A(\U1/aes_core/SB1/n2494 ), .Y(
        \U1/aes_core/SB1/n2444 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1024  ( .A(\U1/aes_core/SB1/n2444 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2234 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1023  ( .AN(\U1/aes_core/SB1/n2207 ), 
        .B(\U1/aes_core/SB1/n2091 ), .C(\U1/aes_core/SB1/n2090 ), .D(
        \U1/aes_core/SB1/n2234 ), .Y(\U1/aes_core/SB1/n2100 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1022  ( .A(\U1/aes_core/SB1/n2103 ), .B(
        \U1/aes_core/SB1/n2101 ), .Y(\U1/aes_core/SB1/n2514 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1021  ( .A(\U1/aes_core/SB1/n2093 ), .B(
        \U1/aes_core/SB1/n2092 ), .Y(\U1/aes_core/SB1/n2506 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U1020  ( .A0(\U1/aes_core/SB1/n2156 ), 
        .A1(\U1/aes_core/SB1/n2308 ), .B0(\U1/aes_core/SB1/n2514 ), .B1(
        \U1/aes_core/SB1/n2423 ), .C0(\U1/aes_core/SB1/n2506 ), .C1(
        \U1/aes_core/SB1/n2441 ), .Y(\U1/aes_core/SB1/n2099 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1019  ( .A(\U1/aes_core/SB1/n2465 ), .B(
        \U1/aes_core/SB1/n2156 ), .Y(\U1/aes_core/SB1/n2292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1018  ( .A(\U1/aes_core/SB1/n2214 ), .B(
        \U1/aes_core/SB1/n2403 ), .Y(\U1/aes_core/SB1/n2245 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1017  ( .A(\U1/aes_core/SB1/n2466 ), .B(
        \U1/aes_core/SB1/n2467 ), .Y(\U1/aes_core/SB1/n2265 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1016  ( .A(\U1/aes_core/SB1/n2421 ), .Y(
        \U1/aes_core/SB1/n2495 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1015  ( .A(\U1/aes_core/SB1/n2495 ), .B(
        \U1/aes_core/SB1/n2300 ), .Y(\U1/aes_core/SB1/n2303 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1014  ( .AN(\U1/aes_core/SB1/n2292 ), 
        .B(\U1/aes_core/SB1/n2245 ), .C(\U1/aes_core/SB1/n2265 ), .D(
        \U1/aes_core/SB1/n2303 ), .Y(\U1/aes_core/SB1/n2098 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1013  ( .A(\U1/aes_core/SB1/n2111 ), .B(
        \U1/aes_core/SB1/n2103 ), .Y(\U1/aes_core/SB1/n2215 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1012  ( .A(\U1/aes_core/SB1/n2215 ), .B(
        \U1/aes_core/SB1/n2477 ), .Y(\U1/aes_core/SB1/n2394 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1011  ( .A(\U1/aes_core/SB1/n2095 ), .B(
        \U1/aes_core/SB1/n2094 ), .Y(\U1/aes_core/SB1/n2513 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1010  ( .A(\U1/aes_core/SB1/n2480 ), .B(
        \U1/aes_core/SB1/n2513 ), .Y(\U1/aes_core/SB1/n2359 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1009  ( .A(\U1/aes_core/SB1/n2359 ), .Y(
        \U1/aes_core/SB1/n2096 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1008  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2300 ), .Y(\U1/aes_core/SB1/n2378 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1007  ( .A(\U1/aes_core/SB1/n2513 ), .Y(
        \U1/aes_core/SB1/n2496 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1006  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2496 ), .Y(\U1/aes_core/SB1/n2429 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U1005  ( .AN(\U1/aes_core/SB1/n2394 ), 
        .B(\U1/aes_core/SB1/n2096 ), .C(\U1/aes_core/SB1/n2378 ), .D(
        \U1/aes_core/SB1/n2429 ), .Y(\U1/aes_core/SB1/n2097 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U1004  ( .A(\U1/aes_core/SB1/n2100 ), .B(
        \U1/aes_core/SB1/n2099 ), .C(\U1/aes_core/SB1/n2098 ), .D(
        \U1/aes_core/SB1/n2097 ), .Y(\U1/aes_core/SB1/n2196 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1003  ( .A(\U1/aes_core/SB1/n2420 ), .B(
        \U1/aes_core/SB1/n2215 ), .Y(\U1/aes_core/SB1/n2428 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U1002  ( .A(\U1/aes_core/SB1/n2110 ), .B(
        \U1/aes_core/SB1/n2101 ), .Y(\U1/aes_core/SB1/n2311 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U1001  ( .A(\U1/aes_core/SB1/n2402 ), .B(
        \U1/aes_core/SB1/n2311 ), .Y(\U1/aes_core/SB1/n2282 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U1000  ( .A(\U1/aes_core/SB1/n2514 ), .Y(
        \U1/aes_core/SB1/n2470 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U999  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2451 ), .Y(\U1/aes_core/SB1/n2231 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U998  ( .A0(\U1/aes_core/SB1/n2311 ), 
        .A1(\U1/aes_core/SB1/n2513 ), .B0(\U1/aes_core/SB1/n2231 ), .Y(
        \U1/aes_core/SB1/n2109 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U997  ( .A(\U1/aes_core/SB1/n2351 ), .Y(
        \U1/aes_core/SB1/n2446 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U996  ( .A(\U1/aes_core/SB1/n2446 ), .B(
        \U1/aes_core/SB1/n2469 ), .Y(\U1/aes_core/SB1/n2447 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U995  ( .A(\U1/aes_core/SB1/n2469 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2406 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U994  ( .A(\U1/aes_core/SB1/n2103 ), .B(
        \U1/aes_core/SB1/n2102 ), .Y(\U1/aes_core/SB1/n2476 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U993  ( .A(\U1/aes_core/SB1/n2476 ), .Y(
        \U1/aes_core/SB1/n2226 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U992  ( .A(\U1/aes_core/SB1/n2442 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2250 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U991  ( .A(\U1/aes_core/SB1/n2464 ), .Y(
        \U1/aes_core/SB1/n2445 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U990  ( .A(\U1/aes_core/SB1/n2445 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2314 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U989  ( .A(\U1/aes_core/SB1/n2447 ), .B(
        \U1/aes_core/SB1/n2406 ), .C(\U1/aes_core/SB1/n2250 ), .D(
        \U1/aes_core/SB1/n2314 ), .Y(\U1/aes_core/SB1/n2108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U988  ( .A(\U1/aes_core/SB1/n2466 ), .B(
        \U1/aes_core/SB1/n2444 ), .Y(\U1/aes_core/SB1/n2373 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U987  ( .A(\U1/aes_core/SB1/n2508 ), .B(
        \U1/aes_core/SB1/n2444 ), .Y(\U1/aes_core/SB1/n2364 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U986  ( .A(\U1/aes_core/SB1/n2506 ), .Y(
        \U1/aes_core/SB1/n2499 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U985  ( .A(\U1/aes_core/SB1/n2403 ), .B(
        \U1/aes_core/SB1/n2499 ), .Y(\U1/aes_core/SB1/n2211 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U984  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2442 ), .Y(\U1/aes_core/SB1/n2347 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U983  ( .A(\U1/aes_core/SB1/n2373 ), .B(
        \U1/aes_core/SB1/n2364 ), .C(\U1/aes_core/SB1/n2211 ), .D(
        \U1/aes_core/SB1/n2347 ), .Y(\U1/aes_core/SB1/n2107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U982  ( .A(\U1/aes_core/SB1/n2418 ), .Y(
        \U1/aes_core/SB1/n2387 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U981  ( .A(\U1/aes_core/SB1/n2214 ), .B(
        \U1/aes_core/SB1/n2387 ), .Y(\U1/aes_core/SB1/n2198 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U980  ( .A(\U1/aes_core/SB1/n2105 ), .B(
        \U1/aes_core/SB1/n2104 ), .Y(\U1/aes_core/SB1/n2453 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U979  ( .A(\U1/aes_core/SB1/n2453 ), .Y(
        \U1/aes_core/SB1/n2487 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U978  ( .A(\U1/aes_core/SB1/n2214 ), .B(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2262 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U977  ( .A(\U1/aes_core/SB1/n2402 ), .Y(
        \U1/aes_core/SB1/n2510 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U976  ( .A(\U1/aes_core/SB1/n2510 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2297 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U975  ( .A(\U1/aes_core/SB1/n2443 ), .B(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2471 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U974  ( .A(\U1/aes_core/SB1/n2198 ), .B(
        \U1/aes_core/SB1/n2262 ), .C(\U1/aes_core/SB1/n2297 ), .D(
        \U1/aes_core/SB1/n2471 ), .Y(\U1/aes_core/SB1/n2106 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U973  ( .A(\U1/aes_core/SB1/n2428 ), .B(
        \U1/aes_core/SB1/n2282 ), .C(\U1/aes_core/SB1/n2109 ), .D(
        \U1/aes_core/SB1/n2108 ), .E(\U1/aes_core/SB1/n2107 ), .F(
        \U1/aes_core/SB1/n2106 ), .Y(\U1/aes_core/SB1/n2185 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U972  ( .A(\U1/aes_core/SB1/n2185 ), .Y(
        \U1/aes_core/SB1/n2120 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U971  ( .A(\U1/aes_core/SB1/n2478 ), .B(
        \U1/aes_core/SB1/n2311 ), .Y(\U1/aes_core/SB1/n2208 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U970  ( .A(\U1/aes_core/SB1/n2111 ), .B(
        \U1/aes_core/SB1/n2110 ), .Y(\U1/aes_core/SB1/n2475 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U969  ( .A(\U1/aes_core/SB1/n2475 ), .B(
        \U1/aes_core/SB1/n2351 ), .Y(\U1/aes_core/SB1/n2360 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U968  ( .A(\U1/aes_core/SB1/n2360 ), .Y(
        \U1/aes_core/SB1/n2113 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U967  ( .A(\U1/aes_core/SB1/n2353 ), .Y(
        \U1/aes_core/SB1/n2500 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U966  ( .A0(\U1/aes_core/SB1/n2226 ), 
        .A1(\U1/aes_core/SB1/n2500 ), .B0(\U1/aes_core/SB1/n2487 ), .Y(
        \U1/aes_core/SB1/n2112 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U965  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2387 ), .Y(\U1/aes_core/SB1/n2233 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U964  ( .AN(\U1/aes_core/SB1/n2208 ), 
        .B(\U1/aes_core/SB1/n2113 ), .C(\U1/aes_core/SB1/n2112 ), .D(
        \U1/aes_core/SB1/n2233 ), .Y(\U1/aes_core/SB1/n2117 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U963  ( .A0(\U1/aes_core/SB1/n2464 ), 
        .A1(\U1/aes_core/SB1/n2512 ), .B0(\U1/aes_core/SB1/n2370 ), .B1(
        \U1/aes_core/SB1/n2418 ), .C0(\U1/aes_core/SB1/n2477 ), .C1(
        \U1/aes_core/SB1/n2494 ), .Y(\U1/aes_core/SB1/n2116 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U962  ( .A(\U1/aes_core/SB1/n2512 ), .B(
        \U1/aes_core/SB1/n2515 ), .Y(\U1/aes_core/SB1/n2273 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U961  ( .A(\U1/aes_core/SB1/n2500 ), .B(
        \U1/aes_core/SB1/n2442 ), .Y(\U1/aes_core/SB1/n2431 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U960  ( .A(\U1/aes_core/SB1/n2403 ), .B(
        \U1/aes_core/SB1/n2500 ), .Y(\U1/aes_core/SB1/n2365 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U959  ( .A(\U1/aes_core/SB1/n2387 ), .B(
        \U1/aes_core/SB1/n2467 ), .Y(\U1/aes_core/SB1/n2212 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U958  ( .AN(\U1/aes_core/SB1/n2273 ), 
        .B(\U1/aes_core/SB1/n2431 ), .C(\U1/aes_core/SB1/n2365 ), .D(
        \U1/aes_core/SB1/n2212 ), .Y(\U1/aes_core/SB1/n2115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U957  ( .A(\U1/aes_core/SB1/n2510 ), .B(
        \U1/aes_core/SB1/n2495 ), .Y(\U1/aes_core/SB1/n2285 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U956  ( .A(\U1/aes_core/SB1/n2387 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2377 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U955  ( .A(\U1/aes_core/SB1/n2214 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U954  ( .A(\U1/aes_core/SB1/n2446 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2298 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U953  ( .A(\U1/aes_core/SB1/n2285 ), .B(
        \U1/aes_core/SB1/n2377 ), .C(\U1/aes_core/SB1/n2253 ), .D(
        \U1/aes_core/SB1/n2298 ), .Y(\U1/aes_core/SB1/n2114 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U952  ( .A(\U1/aes_core/SB1/n2117 ), .B(
        \U1/aes_core/SB1/n2116 ), .C(\U1/aes_core/SB1/n2115 ), .D(
        \U1/aes_core/SB1/n2114 ), .Y(\U1/aes_core/SB1/n2118 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U951  ( .A(\U1/aes_core/SB1/n2118 ), .Y(
        \U1/aes_core/SB1/n2492 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U950  ( .A(\U1/aes_core/SB1/n2508 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2119 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U949  ( .AN(\U1/aes_core/SB1/n2196 ), 
        .B(\U1/aes_core/SB1/n2120 ), .C(\U1/aes_core/SB1/n2492 ), .D(
        \U1/aes_core/SB1/n2119 ), .Y(\U1/aes_core/SB1/n2121 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U948  ( .A(\U1/aes_core/SB1/n2246 ), .B(
        \U1/aes_core/SB1/n2368 ), .C(\U1/aes_core/SB1/n2124 ), .D(
        \U1/aes_core/SB1/n2123 ), .E(\U1/aes_core/SB1/n2122 ), .F(
        \U1/aes_core/SB1/n2121 ), .Y(\U1/aes_core/SB1/n2175 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U947  ( .A(\U1/aes_core/SB1/n2493 ), .B(
        \U1/aes_core/SB1/n2156 ), .Y(\U1/aes_core/SB1/n2291 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U946  ( .A(\U1/aes_core/SB1/n2443 ), .B(
        \U1/aes_core/SB1/n2510 ), .Y(\U1/aes_core/SB1/n2367 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U945  ( .A(\U1/aes_core/SB1/n2499 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2244 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U944  ( .A(\U1/aes_core/SB1/n2215 ), .Y(
        \U1/aes_core/SB1/n2488 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U943  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2267 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U942  ( .AN(\U1/aes_core/SB1/n2291 ), 
        .B(\U1/aes_core/SB1/n2367 ), .C(\U1/aes_core/SB1/n2244 ), .D(
        \U1/aes_core/SB1/n2267 ), .Y(\U1/aes_core/SB1/n2131 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U941  ( .A(\U1/aes_core/SB1/n2480 ), .B(
        \U1/aes_core/SB1/n2351 ), .Y(\U1/aes_core/SB1/n2393 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U940  ( .A(\U1/aes_core/SB1/n2403 ), .B(
        \U1/aes_core/SB1/n2469 ), .Y(\U1/aes_core/SB1/n2224 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U939  ( .A0(\U1/aes_core/SB1/n2489 ), 
        .A1(\U1/aes_core/SB1/n2409 ), .B0(\U1/aes_core/SB1/n2214 ), .Y(
        \U1/aes_core/SB1/n2125 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U938  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2316 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U937  ( .AN(\U1/aes_core/SB1/n2393 ), 
        .B(\U1/aes_core/SB1/n2224 ), .C(\U1/aes_core/SB1/n2125 ), .D(
        \U1/aes_core/SB1/n2316 ), .Y(\U1/aes_core/SB1/n2126 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U936  ( .A(\U1/aes_core/SB1/n2126 ), .Y(
        \U1/aes_core/SB1/n2130 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U935  ( .A(\U1/aes_core/SB1/n2370 ), .Y(
        \U1/aes_core/SB1/n2490 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U934  ( .A(\U1/aes_core/SB1/n2515 ), .Y(
        \U1/aes_core/SB1/n2410 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U933  ( .A0(\U1/aes_core/SB1/n2510 ), 
        .A1(\U1/aes_core/SB1/n2444 ), .B0(\U1/aes_core/SB1/n2490 ), .B1(
        \U1/aes_core/SB1/n2300 ), .C0(\U1/aes_core/SB1/n2410 ), .C1(
        \U1/aes_core/SB1/n2488 ), .Y(\U1/aes_core/SB1/n2129 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U932  ( .A0(\U1/aes_core/SB1/n2311 ), 
        .A1(\U1/aes_core/SB1/n2493 ), .B0(\U1/aes_core/SB1/n2513 ), .B1(
        \U1/aes_core/SB1/n2514 ), .Y(\U1/aes_core/SB1/n2127 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U931  ( .A0(\U1/aes_core/SB1/n2387 ), 
        .A1(\U1/aes_core/SB1/n2200 ), .B0(\U1/aes_core/SB1/n2443 ), .B1(
        \U1/aes_core/SB1/n2466 ), .C0(\U1/aes_core/SB1/n2127 ), .Y(
        \U1/aes_core/SB1/n2128 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U930  ( .AN(\U1/aes_core/SB1/n2131 ), 
        .B(\U1/aes_core/SB1/n2130 ), .C(\U1/aes_core/SB1/n2129 ), .D(
        \U1/aes_core/SB1/n2128 ), .Y(\U1/aes_core/SB1/n2194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U929  ( .A(\U1/aes_core/SB1/n2514 ), .B(
        \U1/aes_core/SB1/n2351 ), .Y(\U1/aes_core/SB1/n2209 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U928  ( .A0(\U1/aes_core/SB1/n2421 ), 
        .A1(\U1/aes_core/SB1/n2514 ), .B0(\U1/aes_core/SB1/n2453 ), .Y(
        \U1/aes_core/SB1/n2136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U927  ( .A(\U1/aes_core/SB1/n2453 ), .B(
        \U1/aes_core/SB1/n2441 ), .Y(\U1/aes_core/SB1/n2293 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB1/U926  ( .A0(\U1/aes_core/SB1/n2442 ), .A1(
        \U1/aes_core/SB1/n2200 ), .B0(\U1/aes_core/SB1/n2293 ), .B1(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2135 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U925  ( .A0(\U1/aes_core/SB1/n2475 ), 
        .A1(\U1/aes_core/SB1/n2515 ), .B0(\U1/aes_core/SB1/n2215 ), .B1(
        \U1/aes_core/SB1/n2308 ), .C0(\U1/aes_core/SB1/n2477 ), .C1(
        \U1/aes_core/SB1/n2506 ), .Y(\U1/aes_core/SB1/n2134 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U924  ( .A(\U1/aes_core/SB1/n2311 ), .Y(
        \U1/aes_core/SB1/n2404 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U923  ( .A(\U1/aes_core/SB1/n2508 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2430 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U922  ( .A(\U1/aes_core/SB1/n2403 ), .B(
        \U1/aes_core/SB1/n2200 ), .Y(\U1/aes_core/SB1/n2232 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U921  ( .A(\U1/aes_core/SB1/n2214 ), .B(
        \U1/aes_core/SB1/n2446 ), .Y(\U1/aes_core/SB1/n2252 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U920  ( .A(\U1/aes_core/SB1/n2403 ), .B(
        \U1/aes_core/SB1/n2444 ), .Y(\U1/aes_core/SB1/n2376 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U919  ( .A(\U1/aes_core/SB1/n2430 ), .B(
        \U1/aes_core/SB1/n2232 ), .C(\U1/aes_core/SB1/n2252 ), .D(
        \U1/aes_core/SB1/n2376 ), .Y(\U1/aes_core/SB1/n2133 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U918  ( .A(\U1/aes_core/SB1/n2423 ), .B(
        \U1/aes_core/SB1/n2311 ), .Y(\U1/aes_core/SB1/n2274 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U917  ( .A(\U1/aes_core/SB1/n2409 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2284 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U916  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2300 ), .Y(\U1/aes_core/SB1/n2315 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U915  ( .AN(\U1/aes_core/SB1/n2274 ), 
        .B(\U1/aes_core/SB1/n2284 ), .C(\U1/aes_core/SB1/n2315 ), .Y(
        \U1/aes_core/SB1/n2132 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U914  ( .A(\U1/aes_core/SB1/n2209 ), .B(
        \U1/aes_core/SB1/n2136 ), .C(\U1/aes_core/SB1/n2135 ), .D(
        \U1/aes_core/SB1/n2134 ), .E(\U1/aes_core/SB1/n2133 ), .F(
        \U1/aes_core/SB1/n2132 ), .Y(\U1/aes_core/SB1/n2521 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U913  ( .A0(\U1/aes_core/SB1/n2214 ), 
        .A1(\U1/aes_core/SB1/n2467 ), .B0(\U1/aes_core/SB1/n2498 ), .Y(
        \U1/aes_core/SB1/n2137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U912  ( .A(\U1/aes_core/SB1/n2200 ), .B(
        \U1/aes_core/SB1/n2300 ), .Y(\U1/aes_core/SB1/n2362 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U911  ( .A(\U1/aes_core/SB1/n2442 ), .B(
        \U1/aes_core/SB1/n2490 ), .Y(\U1/aes_core/SB1/n2229 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U910  ( .A(\U1/aes_core/SB1/n2490 ), .B(
        \U1/aes_core/SB1/n2446 ), .Y(\U1/aes_core/SB1/n2280 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U909  ( .A(\U1/aes_core/SB1/n2137 ), .B(
        \U1/aes_core/SB1/n2362 ), .C(\U1/aes_core/SB1/n2229 ), .D(
        \U1/aes_core/SB1/n2280 ), .Y(\U1/aes_core/SB1/n2141 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U908  ( .A0(\U1/aes_core/SB1/n2493 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2215 ), .B1(
        \U1/aes_core/SB1/n2465 ), .C0(\U1/aes_core/SB1/n2494 ), .C1(
        \U1/aes_core/SB1/n2351 ), .Y(\U1/aes_core/SB1/n2140 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U907  ( .A(\U1/aes_core/SB1/n2445 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2261 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U906  ( .A(\U1/aes_core/SB1/n2444 ), .B(
        \U1/aes_core/SB1/n2496 ), .Y(\U1/aes_core/SB1/n2426 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U905  ( .A(\U1/aes_core/SB1/n2444 ), .B(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U904  ( .A(\U1/aes_core/SB1/n2499 ), .B(
        \U1/aes_core/SB1/n2489 ), .Y(\U1/aes_core/SB1/n2210 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U903  ( .A(\U1/aes_core/SB1/n2261 ), .B(
        \U1/aes_core/SB1/n2426 ), .C(\U1/aes_core/SB1/n2248 ), .D(
        \U1/aes_core/SB1/n2210 ), .Y(\U1/aes_core/SB1/n2139 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U902  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2348 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U901  ( .A(\U1/aes_core/SB1/n2508 ), .B(
        \U1/aes_core/SB1/n2469 ), .Y(\U1/aes_core/SB1/n2296 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U900  ( .A(\U1/aes_core/SB1/n2498 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2372 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U899  ( .A(\U1/aes_core/SB1/n2226 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2197 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U898  ( .A(\U1/aes_core/SB1/n2348 ), .B(
        \U1/aes_core/SB1/n2296 ), .C(\U1/aes_core/SB1/n2372 ), .D(
        \U1/aes_core/SB1/n2197 ), .Y(\U1/aes_core/SB1/n2138 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U897  ( .A(\U1/aes_core/SB1/n2141 ), .B(
        \U1/aes_core/SB1/n2140 ), .C(\U1/aes_core/SB1/n2139 ), .D(
        \U1/aes_core/SB1/n2138 ), .Y(\U1/aes_core/SB1/n2183 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U896  ( .A(\U1/aes_core/SB1/n2175 ), .B(
        \U1/aes_core/SB1/n2194 ), .C(\U1/aes_core/SB1/n2521 ), .D(
        \U1/aes_core/SB1/n2183 ), .Y(\U1/aes_core/SB1/n2150 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U895  ( .A(\U1/aes_core/SB1/n2475 ), .Y(
        \U1/aes_core/SB1/n2399 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U894  ( .A0(\U1/aes_core/SB1/n2351 ), 
        .A1(\U1/aes_core/SB1/n2157 ), .B0(\U1/aes_core/SB1/n2295 ), .B1(
        \U1/aes_core/SB1/n2506 ), .Y(\U1/aes_core/SB1/n2142 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U893  ( .A0(\U1/aes_core/SB1/n2399 ), 
        .A1(\U1/aes_core/SB1/n2451 ), .B0(\U1/aes_core/SB1/n2500 ), .B1(
        \U1/aes_core/SB1/n2508 ), .C0(\U1/aes_core/SB1/n2142 ), .Y(
        \U1/aes_core/SB1/n2149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U892  ( .A(\U1/aes_core/SB1/n2420 ), .B(
        \U1/aes_core/SB1/n2423 ), .Y(\U1/aes_core/SB1/n2419 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U891  ( .A0(\U1/aes_core/SB1/n2354 ), 
        .A1(\U1/aes_core/SB1/n2423 ), .B0(\U1/aes_core/SB1/n2311 ), .B1(
        \U1/aes_core/SB1/n2464 ), .Y(\U1/aes_core/SB1/n2143 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U890  ( .A0(\U1/aes_core/SB1/n2226 ), 
        .A1(\U1/aes_core/SB1/n2419 ), .B0(\U1/aes_core/SB1/n2470 ), .B1(
        \U1/aes_core/SB1/n2489 ), .C0(\U1/aes_core/SB1/n2143 ), .Y(
        \U1/aes_core/SB1/n2148 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U889  ( .A(\U1/aes_core/SB1/n2494 ), .B(
        \U1/aes_core/SB1/n2353 ), .Y(\U1/aes_core/SB1/n2146 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U888  ( .A(\U1/aes_core/SB1/n2444 ), .B(
        \U1/aes_core/SB1/n2469 ), .Y(\U1/aes_core/SB1/n2411 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U887  ( .A(\U1/aes_core/SB1/n2411 ), .Y(
        \U1/aes_core/SB1/n2145 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U886  ( .A(\U1/aes_core/SB1/n2402 ), .B(
        \U1/aes_core/SB1/n2475 ), .Y(\U1/aes_core/SB1/n2258 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U885  ( .A(\U1/aes_core/SB1/n2480 ), .B(
        \U1/aes_core/SB1/n2478 ), .Y(\U1/aes_core/SB1/n2436 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U883  ( .A(\U1/aes_core/SB1/n2451 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2268 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U881  ( .A0(\U1/aes_core/SB1/n2410 ), 
        .A1(\U1/aes_core/SB1/n2146 ), .B0(\U1/aes_core/SB1/n2387 ), .B1(
        \U1/aes_core/SB1/n2145 ), .C0(\U1/aes_core/SB1/n2144 ), .Y(
        \U1/aes_core/SB1/n2147 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U880  ( .AN(\U1/aes_core/SB1/n2150 ), 
        .B(\U1/aes_core/SB1/n2149 ), .C(\U1/aes_core/SB1/n2148 ), .D(
        \U1/aes_core/SB1/n2147 ), .Y(\U1/aes_core/sb1 [16]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U879  ( .A(\U1/aes_core/SB1/n2423 ), .B(
        \U1/aes_core/SB1/n2215 ), .Y(\U1/aes_core/SB1/n2275 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U878  ( .A(\U1/aes_core/SB1/n2370 ), .B(
        \U1/aes_core/SB1/n2420 ), .Y(\U1/aes_core/SB1/n2235 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U877  ( .A(\U1/aes_core/SB1/n2387 ), .B(
        \U1/aes_core/SB1/n2498 ), .Y(\U1/aes_core/SB1/n2369 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U876  ( .A0(\U1/aes_core/SB1/n2369 ), 
        .A1(\U1/aes_core/SB1/n2423 ), .B0(\U1/aes_core/SB1/n2512 ), .Y(
        \U1/aes_core/SB1/n2155 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U875  ( .A(\U1/aes_core/SB1/n2451 ), .B(
        \U1/aes_core/SB1/n2499 ), .Y(\U1/aes_core/SB1/n2251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U874  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2451 ), .Y(\U1/aes_core/SB1/n2375 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U873  ( .A(\U1/aes_core/SB1/n2496 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2283 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U872  ( .A(\U1/aes_core/SB1/n2251 ), .B(
        \U1/aes_core/SB1/n2375 ), .C(\U1/aes_core/SB1/n2283 ), .Y(
        \U1/aes_core/SB1/n2154 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U871  ( .A(\U1/aes_core/SB1/n2451 ), .B(
        \U1/aes_core/SB1/n2510 ), .Y(\U1/aes_core/SB1/n2310 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U870  ( .A(\U1/aes_core/SB1/n2496 ), .B(
        \U1/aes_core/SB1/n2487 ), .C(\U1/aes_core/SB1/n2508 ), .Y(
        \U1/aes_core/SB1/n2151 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U869  ( .A0(\U1/aes_core/SB1/n2310 ), 
        .A1(\U1/aes_core/SB1/n2476 ), .B0(\U1/aes_core/SB1/n2151 ), .B1(
        \U1/aes_core/SB1/n2506 ), .C0(\U1/aes_core/SB1/n2370 ), .C1(
        \U1/aes_core/SB1/n2402 ), .Y(\U1/aes_core/SB1/n2153 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U868  ( .A0(\U1/aes_core/SB1/n2477 ), 
        .A1(\U1/aes_core/SB1/n2505 ), .B0(\U1/aes_core/SB1/n2478 ), .B1(
        \U1/aes_core/SB1/n2475 ), .Y(\U1/aes_core/SB1/n2152 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U867  ( .A(\U1/aes_core/SB1/n2275 ), .B(
        \U1/aes_core/SB1/n2235 ), .C(\U1/aes_core/SB1/n2155 ), .D(
        \U1/aes_core/SB1/n2154 ), .E(\U1/aes_core/SB1/n2153 ), .F(
        \U1/aes_core/SB1/n2152 ), .Y(\U1/aes_core/SB1/n2520 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U866  ( .A(\U1/aes_core/SB1/n2351 ), .B(
        \U1/aes_core/SB1/n2311 ), .Y(\U1/aes_core/SB1/n2201 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U865  ( .A0(\U1/aes_core/SB1/n2351 ), 
        .A1(\U1/aes_core/SB1/n2441 ), .B0(\U1/aes_core/SB1/n2215 ), .Y(
        \U1/aes_core/SB1/n2162 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U864  ( .A(\U1/aes_core/SB1/n2445 ), .B(
        \U1/aes_core/SB1/n2451 ), .Y(\U1/aes_core/SB1/n2203 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U863  ( .A0(\U1/aes_core/SB1/n2308 ), 
        .A1(\U1/aes_core/SB1/n2480 ), .B0(\U1/aes_core/SB1/n2203 ), .B1(
        \U1/aes_core/SB1/n2494 ), .Y(\U1/aes_core/SB1/n2161 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U862  ( .A0(\U1/aes_core/SB1/n2295 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2464 ), .B1(
        \U1/aes_core/SB1/n2370 ), .C0(\U1/aes_core/SB1/n2478 ), .C1(
        \U1/aes_core/SB1/n2421 ), .Y(\U1/aes_core/SB1/n2160 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U861  ( .A(\U1/aes_core/SB1/n2513 ), .B(
        \U1/aes_core/SB1/n2156 ), .Y(\U1/aes_core/SB1/n2259 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U860  ( .A(\U1/aes_core/SB1/n2500 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2266 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U859  ( .A(\U1/aes_core/SB1/n2442 ), .B(
        \U1/aes_core/SB1/n2495 ), .Y(\U1/aes_core/SB1/n2276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U858  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2510 ), .Y(\U1/aes_core/SB1/n2405 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U857  ( .AN(\U1/aes_core/SB1/n2259 ), 
        .B(\U1/aes_core/SB1/n2266 ), .C(\U1/aes_core/SB1/n2276 ), .D(
        \U1/aes_core/SB1/n2405 ), .Y(\U1/aes_core/SB1/n2159 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U856  ( .A(\U1/aes_core/SB1/n2402 ), .B(
        \U1/aes_core/SB1/n2157 ), .Y(\U1/aes_core/SB1/n2384 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U855  ( .A(\U1/aes_core/SB1/n2480 ), .B(
        \U1/aes_core/SB1/n2464 ), .Y(\U1/aes_core/SB1/n2437 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U853  ( .A(\U1/aes_core/SB1/n2200 ), .B(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2225 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U851  ( .A(\U1/aes_core/SB1/n2201 ), .B(
        \U1/aes_core/SB1/n2162 ), .C(\U1/aes_core/SB1/n2161 ), .D(
        \U1/aes_core/SB1/n2160 ), .E(\U1/aes_core/SB1/n2159 ), .F(
        \U1/aes_core/SB1/n2158 ), .Y(\U1/aes_core/SB1/n2195 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U850  ( .A(\U1/aes_core/SB1/n2418 ), .B(
        \U1/aes_core/SB1/n2215 ), .Y(\U1/aes_core/SB1/n2213 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U849  ( .A(\U1/aes_core/SB1/n2370 ), .B(
        \U1/aes_core/SB1/n2295 ), .Y(\U1/aes_core/SB1/n2450 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U848  ( .A(\U1/aes_core/SB1/n2351 ), .B(
        \U1/aes_core/SB1/n2421 ), .Y(\U1/aes_core/SB1/n2263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U847  ( .A(\U1/aes_core/SB1/n2515 ), .B(
        \U1/aes_core/SB1/n2421 ), .Y(\U1/aes_core/SB1/n2278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U846  ( .A(\U1/aes_core/SB1/n2446 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2363 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U845  ( .A(\U1/aes_core/SB1/n2496 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U844  ( .A(\U1/aes_core/SB1/n2500 ), .B(
        \U1/aes_core/SB1/n2496 ), .Y(\U1/aes_core/SB1/n2349 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U843  ( .A(\U1/aes_core/SB1/n2410 ), .B(
        \U1/aes_core/SB1/n2467 ), .Y(\U1/aes_core/SB1/n2249 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U842  ( .A(\U1/aes_core/SB1/n2363 ), .B(
        \U1/aes_core/SB1/n2230 ), .C(\U1/aes_core/SB1/n2349 ), .D(
        \U1/aes_core/SB1/n2249 ), .Y(\U1/aes_core/SB1/n2166 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U841  ( .A(\U1/aes_core/SB1/n2515 ), .B(
        \U1/aes_core/SB1/n2311 ), .Y(\U1/aes_core/SB1/n2299 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U840  ( .A(\U1/aes_core/SB1/n2514 ), .B(
        \U1/aes_core/SB1/n2295 ), .Y(\U1/aes_core/SB1/n2424 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U839  ( .A(\U1/aes_core/SB1/n2441 ), .B(
        \U1/aes_core/SB1/n2480 ), .Y(\U1/aes_core/SB1/n2374 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U838  ( .A(\U1/aes_core/SB1/n2402 ), .B(
        \U1/aes_core/SB1/n2480 ), .Y(\U1/aes_core/SB1/n2199 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U837  ( .A0(\U1/aes_core/SB1/n2480 ), 
        .A1(\U1/aes_core/SB1/n2515 ), .B0(\U1/aes_core/SB1/n2311 ), .B1(
        \U1/aes_core/SB1/n2441 ), .Y(\U1/aes_core/SB1/n2164 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U836  ( .A0(\U1/aes_core/SB1/n2295 ), 
        .A1(\U1/aes_core/SB1/n2512 ), .B0(\U1/aes_core/SB1/n2308 ), .B1(
        \U1/aes_core/SB1/n2370 ), .Y(\U1/aes_core/SB1/n2163 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U835  ( .A(\U1/aes_core/SB1/n2299 ), .B(
        \U1/aes_core/SB1/n2424 ), .C(\U1/aes_core/SB1/n2374 ), .D(
        \U1/aes_core/SB1/n2199 ), .E(\U1/aes_core/SB1/n2164 ), .F(
        \U1/aes_core/SB1/n2163 ), .Y(\U1/aes_core/SB1/n2165 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U834  ( .A(\U1/aes_core/SB1/n2213 ), .B(
        \U1/aes_core/SB1/n2450 ), .C(\U1/aes_core/SB1/n2263 ), .D(
        \U1/aes_core/SB1/n2278 ), .E(\U1/aes_core/SB1/n2166 ), .F(
        \U1/aes_core/SB1/n2165 ), .Y(\U1/aes_core/SB1/n2184 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U833  ( .A0(\U1/aes_core/SB1/n2446 ), 
        .A1(\U1/aes_core/SB1/n2443 ), .B0(\U1/aes_core/SB1/n2499 ), .B1(
        \U1/aes_core/SB1/n2387 ), .C0(\U1/aes_core/SB1/n2184 ), .Y(
        \U1/aes_core/SB1/n2167 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U832  ( .A(\U1/aes_core/SB1/n2167 ), .Y(
        \U1/aes_core/SB1/n2174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U831  ( .A(\U1/aes_core/SB1/n2478 ), .B(
        \U1/aes_core/SB1/n2441 ), .Y(\U1/aes_core/SB1/n2468 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U830  ( .A0(\U1/aes_core/SB1/n2445 ), 
        .A1(\U1/aes_core/SB1/n2468 ), .B0(\U1/aes_core/SB1/n2500 ), .Y(
        \U1/aes_core/SB1/n2170 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U829  ( .A0(\U1/aes_core/SB1/n2410 ), 
        .A1(\U1/aes_core/SB1/n2489 ), .B0(\U1/aes_core/SB1/n2452 ), .Y(
        \U1/aes_core/SB1/n2169 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U828  ( .A0(\U1/aes_core/SB1/n2409 ), 
        .A1(\U1/aes_core/SB1/n2451 ), .B0(\U1/aes_core/SB1/n2495 ), .Y(
        \U1/aes_core/SB1/n2168 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U827  ( .A(\U1/aes_core/SB1/n2442 ), .B(
        \U1/aes_core/SB1/n2488 ), .Y(\U1/aes_core/SB1/n2242 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U826  ( .A(\U1/aes_core/SB1/n2170 ), .B(
        \U1/aes_core/SB1/n2169 ), .C(\U1/aes_core/SB1/n2168 ), .D(
        \U1/aes_core/SB1/n2242 ), .Y(\U1/aes_core/SB1/n2173 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U825  ( .A(\U1/aes_core/SB1/n2487 ), .B(
        \U1/aes_core/SB1/n2403 ), .Y(\U1/aes_core/SB1/n2457 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB1/U824  ( .A(\U1/aes_core/SB1/n2457 ), .B(
        \U1/aes_core/SB1/n2477 ), .C(\U1/aes_core/SB1/n2464 ), .Y(
        \U1/aes_core/SB1/n2171 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U823  ( .A0(\U1/aes_core/SB1/n2441 ), 
        .A1(\U1/aes_core/SB1/n2514 ), .B0(\U1/aes_core/SB1/n2171 ), .B1(
        \U1/aes_core/SB1/n2475 ), .C0(\U1/aes_core/SB1/n2513 ), .C1(
        \U1/aes_core/SB1/n2505 ), .Y(\U1/aes_core/SB1/n2172 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U822  ( .A(\U1/aes_core/SB1/n2520 ), .B(
        \U1/aes_core/SB1/n2195 ), .C(\U1/aes_core/SB1/n2175 ), .D(
        \U1/aes_core/SB1/n2174 ), .E(\U1/aes_core/SB1/n2173 ), .F(
        \U1/aes_core/SB1/n2172 ), .Y(\U1/aes_core/sb1 [17]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U821  ( .A0(\U1/aes_core/SB1/n2469 ), 
        .A1(\U1/aes_core/SB1/n2489 ), .B0(\U1/aes_core/SB1/n2510 ), .B1(
        \U1/aes_core/SB1/n2500 ), .Y(\U1/aes_core/SB1/n2176 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U820  ( .A0(\U1/aes_core/SB1/n2420 ), 
        .A1(\U1/aes_core/SB1/n2514 ), .B0(\U1/aes_core/SB1/n2370 ), .B1(
        \U1/aes_core/SB1/n2441 ), .C0(\U1/aes_core/SB1/n2176 ), .Y(
        \U1/aes_core/SB1/n2182 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U819  ( .A(\U1/aes_core/SB1/n2495 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2279 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U818  ( .A(\U1/aes_core/SB1/n2469 ), .B(
        \U1/aes_core/SB1/n2445 ), .Y(\U1/aes_core/SB1/n2260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U817  ( .A(\U1/aes_core/SB1/n2489 ), .B(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2228 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U816  ( .A(\U1/aes_core/SB1/n2409 ), .B(
        \U1/aes_core/SB1/n2452 ), .Y(\U1/aes_core/SB1/n2247 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U815  ( .A(\U1/aes_core/SB1/n2279 ), .B(
        \U1/aes_core/SB1/n2260 ), .C(\U1/aes_core/SB1/n2228 ), .D(
        \U1/aes_core/SB1/n2247 ), .Y(\U1/aes_core/SB1/n2181 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U814  ( .A(\U1/aes_core/SB1/n2515 ), .B(
        \U1/aes_core/SB1/n2493 ), .Y(\U1/aes_core/SB1/n2398 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U813  ( .A0(\U1/aes_core/SB1/n2446 ), 
        .A1(\U1/aes_core/SB1/n2398 ), .B0(\U1/aes_core/SB1/n2499 ), .Y(
        \U1/aes_core/SB1/n2179 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U812  ( .A0(\U1/aes_core/SB1/n2496 ), 
        .A1(\U1/aes_core/SB1/n2387 ), .B0(\U1/aes_core/SB1/n2399 ), .Y(
        \U1/aes_core/SB1/n2178 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U811  ( .A0(\U1/aes_core/SB1/n2404 ), 
        .A1(\U1/aes_core/SB1/n2444 ), .B0(\U1/aes_core/SB1/n2498 ), .Y(
        \U1/aes_core/SB1/n2177 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U810  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2496 ), .Y(\U1/aes_core/SB1/n2371 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U809  ( .A(\U1/aes_core/SB1/n2179 ), .B(
        \U1/aes_core/SB1/n2178 ), .C(\U1/aes_core/SB1/n2177 ), .D(
        \U1/aes_core/SB1/n2371 ), .Y(\U1/aes_core/SB1/n2180 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U808  ( .A(\U1/aes_core/SB1/n2185 ), .B(
        \U1/aes_core/SB1/n2184 ), .C(\U1/aes_core/SB1/n2183 ), .D(
        \U1/aes_core/SB1/n2182 ), .E(\U1/aes_core/SB1/n2181 ), .F(
        \U1/aes_core/SB1/n2180 ), .Y(\U1/aes_core/SB1/n2519 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U807  ( .A0(\U1/aes_core/SB1/n2300 ), 
        .A1(\U1/aes_core/SB1/n2500 ), .B0(\U1/aes_core/SB1/n2508 ), .B1(
        \U1/aes_core/SB1/n2443 ), .C0(\U1/aes_core/SB1/n2519 ), .Y(
        \U1/aes_core/SB1/n2186 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U806  ( .A(\U1/aes_core/SB1/n2186 ), .Y(
        \U1/aes_core/SB1/n2193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U805  ( .A(\U1/aes_core/SB1/n2452 ), .B(
        \U1/aes_core/SB1/n2214 ), .Y(\U1/aes_core/SB1/n2361 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U804  ( .A1N(\U1/aes_core/SB1/n2361 ), 
        .A0(\U1/aes_core/SB1/n2470 ), .B0(\U1/aes_core/SB1/n2442 ), .Y(
        \U1/aes_core/SB1/n2189 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U803  ( .A0(\U1/aes_core/SB1/n2410 ), 
        .A1(\U1/aes_core/SB1/n2293 ), .B0(\U1/aes_core/SB1/n2469 ), .Y(
        \U1/aes_core/SB1/n2188 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U802  ( .A0(\U1/aes_core/SB1/n2496 ), 
        .A1(\U1/aes_core/SB1/n2451 ), .B0(\U1/aes_core/SB1/n2490 ), .Y(
        \U1/aes_core/SB1/n2187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U801  ( .A(\U1/aes_core/SB1/n2467 ), .B(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2243 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U800  ( .A(\U1/aes_core/SB1/n2189 ), .B(
        \U1/aes_core/SB1/n2188 ), .C(\U1/aes_core/SB1/n2187 ), .D(
        \U1/aes_core/SB1/n2243 ), .Y(\U1/aes_core/SB1/n2192 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U799  ( .A(\U1/aes_core/SB1/n2466 ), .B(
        \U1/aes_core/SB1/n2498 ), .Y(\U1/aes_core/SB1/n2497 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U798  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2444 ), .Y(\U1/aes_core/SB1/n2190 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U797  ( .A0(\U1/aes_core/SB1/n2497 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2190 ), .B1(
        \U1/aes_core/SB1/n2478 ), .C0(\U1/aes_core/SB1/n2421 ), .C1(
        \U1/aes_core/SB1/n2423 ), .Y(\U1/aes_core/SB1/n2191 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U796  ( .A(\U1/aes_core/SB1/n2196 ), .B(
        \U1/aes_core/SB1/n2195 ), .C(\U1/aes_core/SB1/n2194 ), .D(
        \U1/aes_core/SB1/n2193 ), .E(\U1/aes_core/SB1/n2192 ), .F(
        \U1/aes_core/SB1/n2191 ), .Y(\U1/aes_core/sb1 [18]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U795  ( .A(\U1/aes_core/SB1/n2300 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2502 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U794  ( .AN(\U1/aes_core/SB1/n2199 ), 
        .B(\U1/aes_core/SB1/n2198 ), .C(\U1/aes_core/SB1/n2197 ), .D(
        \U1/aes_core/SB1/n2502 ), .Y(\U1/aes_core/SB1/n2206 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U793  ( .A0(\U1/aes_core/SB1/n2200 ), 
        .A1(\U1/aes_core/SB1/n2469 ), .B0(\U1/aes_core/SB1/n2387 ), .Y(
        \U1/aes_core/SB1/n2202 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U790  ( .A(\U1/aes_core/SB1/n2443 ), .B(
        \U1/aes_core/SB1/n2490 ), .Y(\U1/aes_core/SB1/n2454 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U789  ( .A0(\U1/aes_core/SB1/n2308 ), 
        .A1(\U1/aes_core/SB1/n2512 ), .B0(\U1/aes_core/SB1/n2454 ), .B1(
        \U1/aes_core/SB1/n2465 ), .C0(\U1/aes_core/SB1/n2506 ), .C1(
        \U1/aes_core/SB1/n2515 ), .Y(\U1/aes_core/SB1/n2204 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U788  ( .A(\U1/aes_core/SB1/n2209 ), .B(
        \U1/aes_core/SB1/n2208 ), .C(\U1/aes_core/SB1/n2207 ), .D(
        \U1/aes_core/SB1/n2206 ), .E(\U1/aes_core/SB1/n2205 ), .F(
        \U1/aes_core/SB1/n2204 ), .Y(\U1/aes_core/SB1/n2417 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U787  ( .AN(\U1/aes_core/SB1/n2213 ), 
        .B(\U1/aes_core/SB1/n2212 ), .C(\U1/aes_core/SB1/n2211 ), .D(
        \U1/aes_core/SB1/n2210 ), .Y(\U1/aes_core/SB1/n2223 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U786  ( .A0(\U1/aes_core/SB1/n2500 ), 
        .A1(\U1/aes_core/SB1/n2410 ), .B0(\U1/aes_core/SB1/n2495 ), .B1(
        \U1/aes_core/SB1/n2409 ), .C0(\U1/aes_core/SB1/n2214 ), .C1(
        \U1/aes_core/SB1/n2510 ), .Y(\U1/aes_core/SB1/n2222 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U785  ( .A0(\U1/aes_core/SB1/n2464 ), 
        .A1(\U1/aes_core/SB1/n2370 ), .B0(\U1/aes_core/SB1/n2215 ), .B1(
        \U1/aes_core/SB1/n2308 ), .Y(\U1/aes_core/SB1/n2216 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U784  ( .A0(\U1/aes_core/SB1/n2387 ), 
        .A1(\U1/aes_core/SB1/n2404 ), .B0(\U1/aes_core/SB1/n2403 ), .B1(
        \U1/aes_core/SB1/n2467 ), .C0(\U1/aes_core/SB1/n2216 ), .Y(
        \U1/aes_core/SB1/n2221 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U783  ( .A(\U1/aes_core/SB1/n2475 ), .B(
        \U1/aes_core/SB1/n2514 ), .Y(\U1/aes_core/SB1/n2218 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U782  ( .A0(\U1/aes_core/SB1/n2300 ), 
        .A1(\U1/aes_core/SB1/n2219 ), .B0(\U1/aes_core/SB1/n2496 ), .B1(
        \U1/aes_core/SB1/n2218 ), .C0(\U1/aes_core/SB1/n2217 ), .Y(
        \U1/aes_core/SB1/n2220 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U781  ( .AN(\U1/aes_core/SB1/n2223 ), 
        .B(\U1/aes_core/SB1/n2222 ), .C(\U1/aes_core/SB1/n2221 ), .D(
        \U1/aes_core/SB1/n2220 ), .Y(\U1/aes_core/SB1/n2462 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U780  ( .A(\U1/aes_core/SB1/n2224 ), .Y(
        \U1/aes_core/SB1/n2240 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U779  ( .A0(\U1/aes_core/SB1/n2354 ), 
        .A1(\U1/aes_core/SB1/n2423 ), .B0(\U1/aes_core/SB1/n2225 ), .Y(
        \U1/aes_core/SB1/n2239 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U778  ( .A0(\U1/aes_core/SB1/n2496 ), 
        .A1(\U1/aes_core/SB1/n2495 ), .B0(\U1/aes_core/SB1/n2466 ), .B1(
        \U1/aes_core/SB1/n2226 ), .Y(\U1/aes_core/SB1/n2227 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U777  ( .A0(\U1/aes_core/SB1/n2477 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2493 ), .B1(
        \U1/aes_core/SB1/n2505 ), .C0(\U1/aes_core/SB1/n2227 ), .Y(
        \U1/aes_core/SB1/n2238 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U776  ( .A(\U1/aes_core/SB1/n2231 ), .B(
        \U1/aes_core/SB1/n2230 ), .C(\U1/aes_core/SB1/n2229 ), .D(
        \U1/aes_core/SB1/n2228 ), .Y(\U1/aes_core/SB1/n2237 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U775  ( .AN(\U1/aes_core/SB1/n2235 ), 
        .B(\U1/aes_core/SB1/n2234 ), .C(\U1/aes_core/SB1/n2233 ), .D(
        \U1/aes_core/SB1/n2232 ), .Y(\U1/aes_core/SB1/n2236 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U774  ( .A(\U1/aes_core/SB1/n2241 ), .B(
        \U1/aes_core/SB1/n2240 ), .C(\U1/aes_core/SB1/n2239 ), .D(
        \U1/aes_core/SB1/n2238 ), .E(\U1/aes_core/SB1/n2237 ), .F(
        \U1/aes_core/SB1/n2236 ), .Y(\U1/aes_core/SB1/n2366 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U773  ( .A0(\U1/aes_core/SB1/n2453 ), 
        .A1(\U1/aes_core/SB1/n2370 ), .B0(\U1/aes_core/SB1/n2242 ), .Y(
        \U1/aes_core/SB1/n2257 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U772  ( .AN(\U1/aes_core/SB1/n2246 ), 
        .B(\U1/aes_core/SB1/n2245 ), .C(\U1/aes_core/SB1/n2244 ), .D(
        \U1/aes_core/SB1/n2243 ), .Y(\U1/aes_core/SB1/n2256 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U771  ( .A(\U1/aes_core/SB1/n2487 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2501 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U770  ( .A(\U1/aes_core/SB1/n2249 ), .B(
        \U1/aes_core/SB1/n2248 ), .C(\U1/aes_core/SB1/n2247 ), .D(
        \U1/aes_core/SB1/n2501 ), .Y(\U1/aes_core/SB1/n2255 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U769  ( .A(\U1/aes_core/SB1/n2253 ), .B(
        \U1/aes_core/SB1/n2252 ), .C(\U1/aes_core/SB1/n2251 ), .D(
        \U1/aes_core/SB1/n2250 ), .Y(\U1/aes_core/SB1/n2254 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U768  ( .A(\U1/aes_core/SB1/n2259 ), .B(
        \U1/aes_core/SB1/n2258 ), .C(\U1/aes_core/SB1/n2257 ), .D(
        \U1/aes_core/SB1/n2256 ), .E(\U1/aes_core/SB1/n2255 ), .F(
        \U1/aes_core/SB1/n2254 ), .Y(\U1/aes_core/SB1/n2390 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U767  ( .AN(\U1/aes_core/SB1/n2263 ), 
        .B(\U1/aes_core/SB1/n2262 ), .C(\U1/aes_core/SB1/n2261 ), .D(
        \U1/aes_core/SB1/n2260 ), .Y(\U1/aes_core/SB1/n2272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U766  ( .A(\U1/aes_core/SB1/n2267 ), .B(
        \U1/aes_core/SB1/n2266 ), .C(\U1/aes_core/SB1/n2265 ), .D(
        \U1/aes_core/SB1/n2264 ), .Y(\U1/aes_core/SB1/n2271 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U765  ( .A(\U1/aes_core/SB1/n2452 ), .B(
        \U1/aes_core/SB1/n2488 ), .C(\U1/aes_core/SB1/n2490 ), .Y(
        \U1/aes_core/SB1/n2269 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U764  ( .A0(\U1/aes_core/SB1/n2269 ), 
        .A1(\U1/aes_core/SB1/n2478 ), .B0(\U1/aes_core/SB1/n2308 ), .B1(
        \U1/aes_core/SB1/n2514 ), .C0(\U1/aes_core/SB1/n2268 ), .Y(
        \U1/aes_core/SB1/n2270 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U763  ( .A(\U1/aes_core/SB1/n2275 ), .B(
        \U1/aes_core/SB1/n2274 ), .C(\U1/aes_core/SB1/n2273 ), .D(
        \U1/aes_core/SB1/n2272 ), .E(\U1/aes_core/SB1/n2271 ), .F(
        \U1/aes_core/SB1/n2270 ), .Y(\U1/aes_core/SB1/n2438 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U762  ( .A0(\U1/aes_core/SB1/n2308 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2276 ), .Y(
        \U1/aes_core/SB1/n2290 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U761  ( .A0(\U1/aes_core/SB1/n2442 ), 
        .A1(\U1/aes_core/SB1/n2444 ), .B0(\U1/aes_core/SB1/n2499 ), .B1(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U760  ( .A0(\U1/aes_core/SB1/n2353 ), 
        .A1(\U1/aes_core/SB1/n2441 ), .B0(\U1/aes_core/SB1/n2354 ), .B1(
        \U1/aes_core/SB1/n2418 ), .C0(\U1/aes_core/SB1/n2277 ), .Y(
        \U1/aes_core/SB1/n2289 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U759  ( .A(\U1/aes_core/SB1/n2278 ), .Y(
        \U1/aes_core/SB1/n2281 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U758  ( .AN(\U1/aes_core/SB1/n2282 ), 
        .B(\U1/aes_core/SB1/n2281 ), .C(\U1/aes_core/SB1/n2280 ), .D(
        \U1/aes_core/SB1/n2279 ), .Y(\U1/aes_core/SB1/n2288 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U757  ( .A(\U1/aes_core/SB1/n2286 ), .B(
        \U1/aes_core/SB1/n2285 ), .C(\U1/aes_core/SB1/n2284 ), .D(
        \U1/aes_core/SB1/n2283 ), .Y(\U1/aes_core/SB1/n2287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U756  ( .A(\U1/aes_core/SB1/n2292 ), .B(
        \U1/aes_core/SB1/n2291 ), .C(\U1/aes_core/SB1/n2290 ), .D(
        \U1/aes_core/SB1/n2289 ), .E(\U1/aes_core/SB1/n2288 ), .F(
        \U1/aes_core/SB1/n2287 ), .Y(\U1/aes_core/SB1/n2397 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U755  ( .A0(\U1/aes_core/SB1/n2488 ), 
        .A1(\U1/aes_core/SB1/n2293 ), .B0(\U1/aes_core/SB1/n2498 ), .B1(
        \U1/aes_core/SB1/n2444 ), .Y(\U1/aes_core/SB1/n2294 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U754  ( .A0(\U1/aes_core/SB1/n2370 ), 
        .A1(\U1/aes_core/SB1/n2515 ), .B0(\U1/aes_core/SB1/n2295 ), .B1(
        \U1/aes_core/SB1/n2505 ), .C0(\U1/aes_core/SB1/n2294 ), .Y(
        \U1/aes_core/SB1/n2307 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U753  ( .AN(\U1/aes_core/SB1/n2299 ), 
        .B(\U1/aes_core/SB1/n2298 ), .C(\U1/aes_core/SB1/n2297 ), .D(
        \U1/aes_core/SB1/n2296 ), .Y(\U1/aes_core/SB1/n2306 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U752  ( .A0(\U1/aes_core/SB1/n2508 ), 
        .A1(\U1/aes_core/SB1/n2300 ), .B0(\U1/aes_core/SB1/n2499 ), .Y(
        \U1/aes_core/SB1/n2304 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U751  ( .A(\U1/aes_core/SB1/n2475 ), .B(
        \U1/aes_core/SB1/n2480 ), .Y(\U1/aes_core/SB1/n2301 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U750  ( .A0(\U1/aes_core/SB1/n2451 ), 
        .A1(\U1/aes_core/SB1/n2301 ), .B0(\U1/aes_core/SB1/n2452 ), .B1(
        \U1/aes_core/SB1/n2398 ), .Y(\U1/aes_core/SB1/n2302 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U749  ( .A(\U1/aes_core/SB1/n2304 ), .B(
        \U1/aes_core/SB1/n2303 ), .C(\U1/aes_core/SB1/n2302 ), .Y(
        \U1/aes_core/SB1/n2305 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U748  ( .A(\U1/aes_core/SB1/n2390 ), .B(
        \U1/aes_core/SB1/n2438 ), .C(\U1/aes_core/SB1/n2397 ), .D(
        \U1/aes_core/SB1/n2307 ), .E(\U1/aes_core/SB1/n2306 ), .F(
        \U1/aes_core/SB1/n2305 ), .Y(\U1/aes_core/SB1/n2484 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U747  ( .A(\U1/aes_core/SB1/n2417 ), .B(
        \U1/aes_core/SB1/n2462 ), .C(\U1/aes_core/SB1/n2366 ), .D(
        \U1/aes_core/SB1/n2484 ), .Y(\U1/aes_core/SB1/n2321 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U746  ( .A0(\U1/aes_core/SB1/n2464 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2308 ), .B1(
        \U1/aes_core/SB1/n2480 ), .Y(\U1/aes_core/SB1/n2309 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U745  ( .A0(\U1/aes_core/SB1/n2469 ), 
        .A1(\U1/aes_core/SB1/n2487 ), .B0(\U1/aes_core/SB1/n2500 ), .B1(
        \U1/aes_core/SB1/n2508 ), .C0(\U1/aes_core/SB1/n2309 ), .Y(
        \U1/aes_core/SB1/n2320 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U744  ( .A(\U1/aes_core/SB1/n2310 ), .Y(
        \U1/aes_core/SB1/n2313 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U743  ( .A0(\U1/aes_core/SB1/n2311 ), 
        .A1(\U1/aes_core/SB1/n2441 ), .B0(\U1/aes_core/SB1/n2369 ), .B1(
        \U1/aes_core/SB1/n2421 ), .Y(\U1/aes_core/SB1/n2312 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U742  ( .A0(\U1/aes_core/SB1/n2488 ), 
        .A1(\U1/aes_core/SB1/n2313 ), .B0(\U1/aes_core/SB1/n2470 ), .B1(
        \U1/aes_core/SB1/n2419 ), .C0(\U1/aes_core/SB1/n2312 ), .Y(
        \U1/aes_core/SB1/n2319 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U741  ( .A0(\U1/aes_core/SB1/n2510 ), 
        .A1(\U1/aes_core/SB1/n2387 ), .B0(\U1/aes_core/SB1/n2490 ), .Y(
        \U1/aes_core/SB1/n2317 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB1/U740  ( .A(\U1/aes_core/SB1/n2317 ), .B(
        \U1/aes_core/SB1/n2316 ), .C(\U1/aes_core/SB1/n2315 ), .D(
        \U1/aes_core/SB1/n2314 ), .Y(\U1/aes_core/SB1/n2318 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U739  ( .AN(\U1/aes_core/SB1/n2321 ), 
        .B(\U1/aes_core/SB1/n2320 ), .C(\U1/aes_core/SB1/n2319 ), .D(
        \U1/aes_core/SB1/n2318 ), .Y(\U1/aes_core/sb1 [19]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U738  ( .A(\U1/aes_core/SB1/n3166 ), .B(
        \U1/aes_core/SB1/n2983 ), .Y(\U1/aes_core/SB1/n3043 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U737  ( .A(\U1/aes_core/SB1/n3113 ), .B(
        \U1/aes_core/SB1/n3163 ), .Y(\U1/aes_core/SB1/n3003 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U736  ( .A(\U1/aes_core/SB1/n3130 ), .B(
        \U1/aes_core/SB1/n3241 ), .Y(\U1/aes_core/SB1/n3112 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U735  ( .A0(\U1/aes_core/SB1/n3112 ), 
        .A1(\U1/aes_core/SB1/n3166 ), .B0(\U1/aes_core/SB1/n3255 ), .Y(
        \U1/aes_core/SB1/n2326 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U734  ( .A(\U1/aes_core/SB1/n3194 ), .B(
        \U1/aes_core/SB1/n3242 ), .Y(\U1/aes_core/SB1/n3019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U733  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3194 ), .Y(\U1/aes_core/SB1/n3118 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U732  ( .A(\U1/aes_core/SB1/n3239 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3051 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U731  ( .A(\U1/aes_core/SB1/n3019 ), .B(
        \U1/aes_core/SB1/n3118 ), .C(\U1/aes_core/SB1/n3051 ), .Y(
        \U1/aes_core/SB1/n2325 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U730  ( .A(\U1/aes_core/SB1/n3194 ), .B(
        \U1/aes_core/SB1/n3253 ), .Y(\U1/aes_core/SB1/n3078 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U729  ( .A(\U1/aes_core/SB1/n3239 ), .B(
        \U1/aes_core/SB1/n3230 ), .C(\U1/aes_core/SB1/n3251 ), .Y(
        \U1/aes_core/SB1/n2322 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U728  ( .A0(\U1/aes_core/SB1/n3078 ), 
        .A1(\U1/aes_core/SB1/n3219 ), .B0(\U1/aes_core/SB1/n2322 ), .B1(
        \U1/aes_core/SB1/n3249 ), .C0(\U1/aes_core/SB1/n3113 ), .C1(
        \U1/aes_core/SB1/n3145 ), .Y(\U1/aes_core/SB1/n2324 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U727  ( .A0(\U1/aes_core/SB1/n3220 ), 
        .A1(\U1/aes_core/SB1/n3248 ), .B0(\U1/aes_core/SB1/n3221 ), .B1(
        \U1/aes_core/SB1/n3218 ), .Y(\U1/aes_core/SB1/n2323 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U726  ( .A(\U1/aes_core/SB1/n3043 ), .B(
        \U1/aes_core/SB1/n3003 ), .C(\U1/aes_core/SB1/n2326 ), .D(
        \U1/aes_core/SB1/n2325 ), .E(\U1/aes_core/SB1/n2324 ), .F(
        \U1/aes_core/SB1/n2323 ), .Y(\U1/aes_core/SB1/n3263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U725  ( .A(\U1/aes_core/SB1/n3094 ), .B(
        \U1/aes_core/SB1/n3079 ), .Y(\U1/aes_core/SB1/n2969 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U724  ( .A0(\U1/aes_core/SB1/n3094 ), 
        .A1(\U1/aes_core/SB1/n3184 ), .B0(\U1/aes_core/SB1/n2983 ), .Y(
        \U1/aes_core/SB1/n2333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U723  ( .A(\U1/aes_core/SB1/n3188 ), .B(
        \U1/aes_core/SB1/n3194 ), .Y(\U1/aes_core/SB1/n2971 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U722  ( .A0(\U1/aes_core/SB1/n3076 ), 
        .A1(\U1/aes_core/SB1/n3223 ), .B0(\U1/aes_core/SB1/n2971 ), .B1(
        \U1/aes_core/SB1/n3237 ), .Y(\U1/aes_core/SB1/n2332 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U721  ( .A0(\U1/aes_core/SB1/n3063 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3207 ), .B1(
        \U1/aes_core/SB1/n3113 ), .C0(\U1/aes_core/SB1/n3221 ), .C1(
        \U1/aes_core/SB1/n3164 ), .Y(\U1/aes_core/SB1/n2331 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U720  ( .A(\U1/aes_core/SB1/n3256 ), .B(
        \U1/aes_core/SB1/n2327 ), .Y(\U1/aes_core/SB1/n3027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U719  ( .A(\U1/aes_core/SB1/n3243 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U718  ( .A(\U1/aes_core/SB1/n3185 ), .B(
        \U1/aes_core/SB1/n3238 ), .Y(\U1/aes_core/SB1/n3044 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U717  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3253 ), .Y(\U1/aes_core/SB1/n3148 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U716  ( .AN(\U1/aes_core/SB1/n3027 ), 
        .B(\U1/aes_core/SB1/n3034 ), .C(\U1/aes_core/SB1/n3044 ), .D(
        \U1/aes_core/SB1/n3148 ), .Y(\U1/aes_core/SB1/n2330 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U715  ( .A(\U1/aes_core/SB1/n3145 ), .B(
        \U1/aes_core/SB1/n2328 ), .Y(\U1/aes_core/SB1/n3127 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U714  ( .A(\U1/aes_core/SB1/n3223 ), .B(
        \U1/aes_core/SB1/n3207 ), .Y(\U1/aes_core/SB1/n3180 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U712  ( .A(\U1/aes_core/SB1/n2968 ), .B(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n2993 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U710  ( .A(\U1/aes_core/SB1/n2969 ), .B(
        \U1/aes_core/SB1/n2333 ), .C(\U1/aes_core/SB1/n2332 ), .D(
        \U1/aes_core/SB1/n2331 ), .E(\U1/aes_core/SB1/n2330 ), .F(
        \U1/aes_core/SB1/n2329 ), .Y(\U1/aes_core/SB1/n2904 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U709  ( .A(\U1/aes_core/SB1/n3161 ), .B(
        \U1/aes_core/SB1/n2983 ), .Y(\U1/aes_core/SB1/n2981 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U708  ( .A(\U1/aes_core/SB1/n3113 ), .B(
        \U1/aes_core/SB1/n3063 ), .Y(\U1/aes_core/SB1/n3193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U707  ( .A(\U1/aes_core/SB1/n3094 ), .B(
        \U1/aes_core/SB1/n3164 ), .Y(\U1/aes_core/SB1/n3031 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U706  ( .A(\U1/aes_core/SB1/n3258 ), .B(
        \U1/aes_core/SB1/n3164 ), .Y(\U1/aes_core/SB1/n3046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U705  ( .A(\U1/aes_core/SB1/n3189 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n3106 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U704  ( .A(\U1/aes_core/SB1/n3239 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n2998 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U703  ( .A(\U1/aes_core/SB1/n3243 ), .B(
        \U1/aes_core/SB1/n3239 ), .Y(\U1/aes_core/SB1/n3092 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U702  ( .A(\U1/aes_core/SB1/n3153 ), .B(
        \U1/aes_core/SB1/n3210 ), .Y(\U1/aes_core/SB1/n3017 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U701  ( .A(\U1/aes_core/SB1/n3106 ), .B(
        \U1/aes_core/SB1/n2998 ), .C(\U1/aes_core/SB1/n3092 ), .D(
        \U1/aes_core/SB1/n3017 ), .Y(\U1/aes_core/SB1/n2337 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U700  ( .A(\U1/aes_core/SB1/n3258 ), .B(
        \U1/aes_core/SB1/n3079 ), .Y(\U1/aes_core/SB1/n3067 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U699  ( .A(\U1/aes_core/SB1/n3257 ), .B(
        \U1/aes_core/SB1/n3063 ), .Y(\U1/aes_core/SB1/n3167 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U698  ( .A(\U1/aes_core/SB1/n3184 ), .B(
        \U1/aes_core/SB1/n3223 ), .Y(\U1/aes_core/SB1/n3117 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U697  ( .A(\U1/aes_core/SB1/n3145 ), .B(
        \U1/aes_core/SB1/n3223 ), .Y(\U1/aes_core/SB1/n2967 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U696  ( .A0(\U1/aes_core/SB1/n3223 ), 
        .A1(\U1/aes_core/SB1/n3258 ), .B0(\U1/aes_core/SB1/n3079 ), .B1(
        \U1/aes_core/SB1/n3184 ), .Y(\U1/aes_core/SB1/n2335 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U695  ( .A0(\U1/aes_core/SB1/n3063 ), 
        .A1(\U1/aes_core/SB1/n3255 ), .B0(\U1/aes_core/SB1/n3076 ), .B1(
        \U1/aes_core/SB1/n3113 ), .Y(\U1/aes_core/SB1/n2334 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U694  ( .A(\U1/aes_core/SB1/n3067 ), .B(
        \U1/aes_core/SB1/n3167 ), .C(\U1/aes_core/SB1/n3117 ), .D(
        \U1/aes_core/SB1/n2967 ), .E(\U1/aes_core/SB1/n2335 ), .F(
        \U1/aes_core/SB1/n2334 ), .Y(\U1/aes_core/SB1/n2336 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U693  ( .A(\U1/aes_core/SB1/n2981 ), .B(
        \U1/aes_core/SB1/n3193 ), .C(\U1/aes_core/SB1/n3031 ), .D(
        \U1/aes_core/SB1/n3046 ), .E(\U1/aes_core/SB1/n2337 ), .F(
        \U1/aes_core/SB1/n2336 ), .Y(\U1/aes_core/SB1/n2893 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U692  ( .A0(\U1/aes_core/SB1/n3189 ), 
        .A1(\U1/aes_core/SB1/n3186 ), .B0(\U1/aes_core/SB1/n3242 ), .B1(
        \U1/aes_core/SB1/n3130 ), .C0(\U1/aes_core/SB1/n2893 ), .Y(
        \U1/aes_core/SB1/n2338 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U691  ( .A(\U1/aes_core/SB1/n2338 ), .Y(
        \U1/aes_core/SB1/n2345 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U690  ( .A(\U1/aes_core/SB1/n3221 ), .B(
        \U1/aes_core/SB1/n3184 ), .Y(\U1/aes_core/SB1/n3211 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U689  ( .A0(\U1/aes_core/SB1/n3188 ), 
        .A1(\U1/aes_core/SB1/n3211 ), .B0(\U1/aes_core/SB1/n3243 ), .Y(
        \U1/aes_core/SB1/n2341 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U688  ( .A0(\U1/aes_core/SB1/n3153 ), 
        .A1(\U1/aes_core/SB1/n3232 ), .B0(\U1/aes_core/SB1/n3195 ), .Y(
        \U1/aes_core/SB1/n2340 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U687  ( .A0(\U1/aes_core/SB1/n3152 ), 
        .A1(\U1/aes_core/SB1/n3194 ), .B0(\U1/aes_core/SB1/n3238 ), .Y(
        \U1/aes_core/SB1/n2339 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U686  ( .A(\U1/aes_core/SB1/n3185 ), .B(
        \U1/aes_core/SB1/n3231 ), .Y(\U1/aes_core/SB1/n3010 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U685  ( .A(\U1/aes_core/SB1/n2341 ), .B(
        \U1/aes_core/SB1/n2340 ), .C(\U1/aes_core/SB1/n2339 ), .D(
        \U1/aes_core/SB1/n3010 ), .Y(\U1/aes_core/SB1/n2344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U684  ( .A(\U1/aes_core/SB1/n3230 ), .B(
        \U1/aes_core/SB1/n3146 ), .Y(\U1/aes_core/SB1/n3200 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB1/U683  ( .A(\U1/aes_core/SB1/n3200 ), .B(
        \U1/aes_core/SB1/n3220 ), .C(\U1/aes_core/SB1/n3207 ), .Y(
        \U1/aes_core/SB1/n2342 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U682  ( .A0(\U1/aes_core/SB1/n3184 ), 
        .A1(\U1/aes_core/SB1/n3257 ), .B0(\U1/aes_core/SB1/n2342 ), .B1(
        \U1/aes_core/SB1/n3218 ), .C0(\U1/aes_core/SB1/n3256 ), .C1(
        \U1/aes_core/SB1/n3248 ), .Y(\U1/aes_core/SB1/n2343 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U681  ( .A(\U1/aes_core/SB1/n3263 ), .B(
        \U1/aes_core/SB1/n2904 ), .C(\U1/aes_core/SB1/n2346 ), .D(
        \U1/aes_core/SB1/n2345 ), .E(\U1/aes_core/SB1/n2344 ), .F(
        \U1/aes_core/SB1/n2343 ), .Y(\U1/aes_core/sb1 [1]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U680  ( .A0(\U1/aes_core/SB1/n2361 ), 
        .A1(\U1/aes_core/SB1/n2476 ), .B0(\U1/aes_core/SB1/n2420 ), .Y(
        \U1/aes_core/SB1/n2358 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U679  ( .A(\U1/aes_core/SB1/n2349 ), .B(
        \U1/aes_core/SB1/n2348 ), .C(\U1/aes_core/SB1/n2347 ), .Y(
        \U1/aes_core/SB1/n2357 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U678  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2499 ), .Y(\U1/aes_core/SB1/n2352 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U677  ( .A(\U1/aes_core/SB1/n2470 ), .B(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2350 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U676  ( .A0(\U1/aes_core/SB1/n2352 ), 
        .A1(\U1/aes_core/SB1/n2351 ), .B0(\U1/aes_core/SB1/n2350 ), .B1(
        \U1/aes_core/SB1/n2493 ), .C0(\U1/aes_core/SB1/n2476 ), .C1(
        \U1/aes_core/SB1/n2402 ), .Y(\U1/aes_core/SB1/n2356 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U675  ( .A0(\U1/aes_core/SB1/n2453 ), 
        .A1(\U1/aes_core/SB1/n2354 ), .B0(\U1/aes_core/SB1/n2515 ), .B1(
        \U1/aes_core/SB1/n2505 ), .C0(\U1/aes_core/SB1/n2478 ), .C1(
        \U1/aes_core/SB1/n2353 ), .Y(\U1/aes_core/SB1/n2355 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U674  ( .A(\U1/aes_core/SB1/n2360 ), .B(
        \U1/aes_core/SB1/n2359 ), .C(\U1/aes_core/SB1/n2358 ), .D(
        \U1/aes_core/SB1/n2357 ), .E(\U1/aes_core/SB1/n2356 ), .F(
        \U1/aes_core/SB1/n2355 ), .Y(\U1/aes_core/SB1/n2485 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U673  ( .A0(\U1/aes_core/SB1/n2361 ), 
        .A1(\U1/aes_core/SB1/n2370 ), .B0(\U1/aes_core/SB1/n2441 ), .Y(
        \U1/aes_core/SB1/n2396 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB1/U672  ( .A0(\U1/aes_core/SB1/n2465 ), 
        .A1(\U1/aes_core/SB1/n2478 ), .A2(\U1/aes_core/SB1/n2418 ), .B0(
        \U1/aes_core/SB1/n2494 ), .Y(\U1/aes_core/SB1/n2395 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U671  ( .A(\U1/aes_core/SB1/n2365 ), .B(
        \U1/aes_core/SB1/n2364 ), .C(\U1/aes_core/SB1/n2363 ), .D(
        \U1/aes_core/SB1/n2362 ), .Y(\U1/aes_core/SB1/n2392 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U670  ( .A(\U1/aes_core/SB1/n2366 ), .Y(
        \U1/aes_core/SB1/n2389 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U669  ( .A(\U1/aes_core/SB1/n2367 ), .Y(
        \U1/aes_core/SB1/n2383 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB1/U668  ( .A0(\U1/aes_core/SB1/n2369 ), 
        .A1(\U1/aes_core/SB1/n2506 ), .B0N(\U1/aes_core/SB1/n2368 ), .Y(
        \U1/aes_core/SB1/n2382 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U667  ( .A0(\U1/aes_core/SB1/n2513 ), 
        .A1(\U1/aes_core/SB1/n2370 ), .B0(\U1/aes_core/SB1/n2420 ), .B1(
        \U1/aes_core/SB1/n2480 ), .C0(\U1/aes_core/SB1/n2494 ), .C1(
        \U1/aes_core/SB1/n2515 ), .Y(\U1/aes_core/SB1/n2381 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U666  ( .AN(\U1/aes_core/SB1/n2374 ), 
        .B(\U1/aes_core/SB1/n2373 ), .C(\U1/aes_core/SB1/n2372 ), .D(
        \U1/aes_core/SB1/n2371 ), .Y(\U1/aes_core/SB1/n2380 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U665  ( .A(\U1/aes_core/SB1/n2378 ), .B(
        \U1/aes_core/SB1/n2377 ), .C(\U1/aes_core/SB1/n2376 ), .D(
        \U1/aes_core/SB1/n2375 ), .Y(\U1/aes_core/SB1/n2379 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U664  ( .A(\U1/aes_core/SB1/n2384 ), .B(
        \U1/aes_core/SB1/n2383 ), .C(\U1/aes_core/SB1/n2382 ), .D(
        \U1/aes_core/SB1/n2381 ), .E(\U1/aes_core/SB1/n2380 ), .F(
        \U1/aes_core/SB1/n2379 ), .Y(\U1/aes_core/SB1/n2385 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U663  ( .A(\U1/aes_core/SB1/n2385 ), .Y(
        \U1/aes_core/SB1/n2463 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U662  ( .A0(\U1/aes_core/SB1/n2453 ), 
        .A1(\U1/aes_core/SB1/n2475 ), .B0(\U1/aes_core/SB1/n2515 ), .B1(
        \U1/aes_core/SB1/n2514 ), .Y(\U1/aes_core/SB1/n2386 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U661  ( .A0(\U1/aes_core/SB1/n2443 ), 
        .A1(\U1/aes_core/SB1/n2387 ), .B0(\U1/aes_core/SB1/n2467 ), .B1(
        \U1/aes_core/SB1/n2489 ), .C0(\U1/aes_core/SB1/n2386 ), .Y(
        \U1/aes_core/SB1/n2388 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U660  ( .AN(\U1/aes_core/SB1/n2390 ), 
        .B(\U1/aes_core/SB1/n2389 ), .C(\U1/aes_core/SB1/n2463 ), .D(
        \U1/aes_core/SB1/n2388 ), .Y(\U1/aes_core/SB1/n2391 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U659  ( .A(\U1/aes_core/SB1/n2396 ), .B(
        \U1/aes_core/SB1/n2395 ), .C(\U1/aes_core/SB1/n2394 ), .D(
        \U1/aes_core/SB1/n2393 ), .E(\U1/aes_core/SB1/n2392 ), .F(
        \U1/aes_core/SB1/n2391 ), .Y(\U1/aes_core/SB1/n2461 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U658  ( .A(\U1/aes_core/SB1/n2397 ), .Y(
        \U1/aes_core/SB1/n2401 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U657  ( .A0(\U1/aes_core/SB1/n2399 ), 
        .A1(\U1/aes_core/SB1/n2398 ), .B0(\U1/aes_core/SB1/n2445 ), .B1(
        \U1/aes_core/SB1/n2404 ), .Y(\U1/aes_core/SB1/n2400 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U656  ( .A0(\U1/aes_core/SB1/n2494 ), 
        .A1(\U1/aes_core/SB1/n2402 ), .B0(\U1/aes_core/SB1/n2401 ), .C0(
        \U1/aes_core/SB1/n2400 ), .Y(\U1/aes_core/SB1/n2416 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U655  ( .A0(\U1/aes_core/SB1/n2403 ), 
        .A1(\U1/aes_core/SB1/n2466 ), .B0(\U1/aes_core/SB1/n2495 ), .Y(
        \U1/aes_core/SB1/n2408 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U654  ( .A0(\U1/aes_core/SB1/n2404 ), 
        .A1(\U1/aes_core/SB1/n2469 ), .B0(\U1/aes_core/SB1/n2498 ), .Y(
        \U1/aes_core/SB1/n2407 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U653  ( .A(\U1/aes_core/SB1/n2408 ), .B(
        \U1/aes_core/SB1/n2407 ), .C(\U1/aes_core/SB1/n2406 ), .D(
        \U1/aes_core/SB1/n2405 ), .Y(\U1/aes_core/SB1/n2415 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U652  ( .A(\U1/aes_core/SB1/n2446 ), .B(
        \U1/aes_core/SB1/n2409 ), .Y(\U1/aes_core/SB1/n2413 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U651  ( .A(\U1/aes_core/SB1/n2410 ), .B(
        \U1/aes_core/SB1/n2451 ), .Y(\U1/aes_core/SB1/n2412 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U650  ( .A0(\U1/aes_core/SB1/n2413 ), 
        .A1(\U1/aes_core/SB1/n2512 ), .B0(\U1/aes_core/SB1/n2412 ), .B1(
        \U1/aes_core/SB1/n2476 ), .C0(\U1/aes_core/SB1/n2411 ), .C1(
        \U1/aes_core/SB1/n2477 ), .Y(\U1/aes_core/SB1/n2414 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U649  ( .A(\U1/aes_core/SB1/n2485 ), .B(
        \U1/aes_core/SB1/n2461 ), .C(\U1/aes_core/SB1/n2417 ), .D(
        \U1/aes_core/SB1/n2416 ), .E(\U1/aes_core/SB1/n2415 ), .F(
        \U1/aes_core/SB1/n2414 ), .Y(\U1/aes_core/sb1 [20]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U648  ( .A1N(\U1/aes_core/SB1/n2419 ), 
        .A0(\U1/aes_core/SB1/n2418 ), .B0(\U1/aes_core/SB1/n2475 ), .Y(
        \U1/aes_core/SB1/n2435 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U647  ( .A(\U1/aes_core/SB1/n2488 ), .B(
        \U1/aes_core/SB1/n2469 ), .Y(\U1/aes_core/SB1/n2422 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U646  ( .A0(\U1/aes_core/SB1/n2512 ), 
        .A1(\U1/aes_core/SB1/n2423 ), .B0(\U1/aes_core/SB1/n2422 ), .B1(
        \U1/aes_core/SB1/n2515 ), .C0(\U1/aes_core/SB1/n2421 ), .C1(
        \U1/aes_core/SB1/n2420 ), .Y(\U1/aes_core/SB1/n2434 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U645  ( .A(\U1/aes_core/SB1/n2424 ), .Y(
        \U1/aes_core/SB1/n2427 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U644  ( .AN(\U1/aes_core/SB1/n2428 ), 
        .B(\U1/aes_core/SB1/n2427 ), .C(\U1/aes_core/SB1/n2426 ), .D(
        \U1/aes_core/SB1/n2425 ), .Y(\U1/aes_core/SB1/n2433 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U643  ( .A(\U1/aes_core/SB1/n2431 ), .B(
        \U1/aes_core/SB1/n2430 ), .C(\U1/aes_core/SB1/n2429 ), .Y(
        \U1/aes_core/SB1/n2432 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U642  ( .A(\U1/aes_core/SB1/n2437 ), .B(
        \U1/aes_core/SB1/n2436 ), .C(\U1/aes_core/SB1/n2435 ), .D(
        \U1/aes_core/SB1/n2434 ), .E(\U1/aes_core/SB1/n2433 ), .F(
        \U1/aes_core/SB1/n2432 ), .Y(\U1/aes_core/SB1/n2486 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U641  ( .A(\U1/aes_core/SB1/n2438 ), .Y(
        \U1/aes_core/SB1/n2440 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U640  ( .A0(\U1/aes_core/SB1/n2499 ), 
        .A1(\U1/aes_core/SB1/n2496 ), .B0(\U1/aes_core/SB1/n2500 ), .B1(
        \U1/aes_core/SB1/n2498 ), .Y(\U1/aes_core/SB1/n2439 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U639  ( .A0(\U1/aes_core/SB1/n2475 ), 
        .A1(\U1/aes_core/SB1/n2441 ), .B0(\U1/aes_core/SB1/n2440 ), .C0(
        \U1/aes_core/SB1/n2439 ), .Y(\U1/aes_core/SB1/n2460 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U638  ( .A0(\U1/aes_core/SB1/n2443 ), 
        .A1(\U1/aes_core/SB1/n2499 ), .B0(\U1/aes_core/SB1/n2442 ), .Y(
        \U1/aes_core/SB1/n2449 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U637  ( .A0(\U1/aes_core/SB1/n2446 ), 
        .A1(\U1/aes_core/SB1/n2445 ), .B0(\U1/aes_core/SB1/n2444 ), .Y(
        \U1/aes_core/SB1/n2448 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U636  ( .AN(\U1/aes_core/SB1/n2450 ), 
        .B(\U1/aes_core/SB1/n2449 ), .C(\U1/aes_core/SB1/n2448 ), .D(
        \U1/aes_core/SB1/n2447 ), .Y(\U1/aes_core/SB1/n2459 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U635  ( .A0(\U1/aes_core/SB1/n2495 ), 
        .A1(\U1/aes_core/SB1/n2452 ), .B0(\U1/aes_core/SB1/n2451 ), .Y(
        \U1/aes_core/SB1/n2456 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB1/U634  ( .A0(\U1/aes_core/SB1/n2477 ), .A1(
        \U1/aes_core/SB1/n2454 ), .B0(\U1/aes_core/SB1/n2514 ), .B1(
        \U1/aes_core/SB1/n2453 ), .Y(\U1/aes_core/SB1/n2455 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U633  ( .A0(\U1/aes_core/SB1/n2457 ), 
        .A1(\U1/aes_core/SB1/n2476 ), .B0(\U1/aes_core/SB1/n2456 ), .C0(
        \U1/aes_core/SB1/n2455 ), .Y(\U1/aes_core/SB1/n2458 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U632  ( .A(\U1/aes_core/SB1/n2486 ), .B(
        \U1/aes_core/SB1/n2462 ), .C(\U1/aes_core/SB1/n2461 ), .D(
        \U1/aes_core/SB1/n2460 ), .E(\U1/aes_core/SB1/n2459 ), .F(
        \U1/aes_core/SB1/n2458 ), .Y(\U1/aes_core/sb1 [21]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U631  ( .A0(\U1/aes_core/SB1/n2465 ), 
        .A1(\U1/aes_core/SB1/n2505 ), .B0(\U1/aes_core/SB1/n2464 ), .B1(
        \U1/aes_core/SB1/n2512 ), .C0(\U1/aes_core/SB1/n2463 ), .Y(
        \U1/aes_core/SB1/n2483 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U630  ( .A0(\U1/aes_core/SB1/n2466 ), 
        .A1(\U1/aes_core/SB1/n2510 ), .B0(\U1/aes_core/SB1/n2499 ), .Y(
        \U1/aes_core/SB1/n2474 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U629  ( .A0(\U1/aes_core/SB1/n2490 ), 
        .A1(\U1/aes_core/SB1/n2467 ), .B0(\U1/aes_core/SB1/n2498 ), .Y(
        \U1/aes_core/SB1/n2473 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U628  ( .A0(\U1/aes_core/SB1/n2470 ), 
        .A1(\U1/aes_core/SB1/n2469 ), .B0(\U1/aes_core/SB1/n2468 ), .Y(
        \U1/aes_core/SB1/n2472 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U627  ( .A(\U1/aes_core/SB1/n2474 ), .B(
        \U1/aes_core/SB1/n2473 ), .C(\U1/aes_core/SB1/n2472 ), .D(
        \U1/aes_core/SB1/n2471 ), .Y(\U1/aes_core/SB1/n2482 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U626  ( .A(\U1/aes_core/SB1/n2505 ), .B(
        \U1/aes_core/SB1/n2475 ), .Y(\U1/aes_core/SB1/n2507 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U625  ( .A(\U1/aes_core/SB1/n2495 ), .B(
        \U1/aes_core/SB1/n2507 ), .Y(\U1/aes_core/SB1/n2479 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U624  ( .A0(\U1/aes_core/SB1/n2493 ), 
        .A1(\U1/aes_core/SB1/n2480 ), .B0(\U1/aes_core/SB1/n2479 ), .B1(
        \U1/aes_core/SB1/n2478 ), .C0(\U1/aes_core/SB1/n2477 ), .C1(
        \U1/aes_core/SB1/n2476 ), .Y(\U1/aes_core/SB1/n2481 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U623  ( .A(\U1/aes_core/SB1/n2486 ), .B(
        \U1/aes_core/SB1/n2485 ), .C(\U1/aes_core/SB1/n2484 ), .D(
        \U1/aes_core/SB1/n2483 ), .E(\U1/aes_core/SB1/n2482 ), .F(
        \U1/aes_core/SB1/n2481 ), .Y(\U1/aes_core/sb1 [22]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U622  ( .A0(\U1/aes_core/SB1/n2490 ), 
        .A1(\U1/aes_core/SB1/n2489 ), .B0(\U1/aes_core/SB1/n2488 ), .B1(
        \U1/aes_core/SB1/n2487 ), .Y(\U1/aes_core/SB1/n2491 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U621  ( .A0(\U1/aes_core/SB1/n2494 ), 
        .A1(\U1/aes_core/SB1/n2493 ), .B0(\U1/aes_core/SB1/n2492 ), .C0(
        \U1/aes_core/SB1/n2491 ), .Y(\U1/aes_core/SB1/n2518 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U620  ( .A1N(\U1/aes_core/SB1/n2497 ), 
        .A0(\U1/aes_core/SB1/n2496 ), .B0(\U1/aes_core/SB1/n2495 ), .Y(
        \U1/aes_core/SB1/n2504 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U619  ( .A0(\U1/aes_core/SB1/n2500 ), 
        .A1(\U1/aes_core/SB1/n2499 ), .B0(\U1/aes_core/SB1/n2498 ), .Y(
        \U1/aes_core/SB1/n2503 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U618  ( .A(\U1/aes_core/SB1/n2504 ), .B(
        \U1/aes_core/SB1/n2503 ), .C(\U1/aes_core/SB1/n2502 ), .D(
        \U1/aes_core/SB1/n2501 ), .Y(\U1/aes_core/SB1/n2517 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U617  ( .A(\U1/aes_core/SB1/n2506 ), .B(
        \U1/aes_core/SB1/n2505 ), .Y(\U1/aes_core/SB1/n2509 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U616  ( .A0(\U1/aes_core/SB1/n2510 ), 
        .A1(\U1/aes_core/SB1/n2509 ), .B0(\U1/aes_core/SB1/n2508 ), .B1(
        \U1/aes_core/SB1/n2507 ), .Y(\U1/aes_core/SB1/n2511 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U615  ( .A0(\U1/aes_core/SB1/n2515 ), 
        .A1(\U1/aes_core/SB1/n2514 ), .B0(\U1/aes_core/SB1/n2513 ), .B1(
        \U1/aes_core/SB1/n2512 ), .C0(\U1/aes_core/SB1/n2511 ), .Y(
        \U1/aes_core/SB1/n2516 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U614  ( .A(\U1/aes_core/SB1/n2521 ), .B(
        \U1/aes_core/SB1/n2520 ), .C(\U1/aes_core/SB1/n2519 ), .D(
        \U1/aes_core/SB1/n2518 ), .E(\U1/aes_core/SB1/n2517 ), .F(
        \U1/aes_core/SB1/n2516 ), .Y(\U1/aes_core/sb1 [23]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U613  ( .A(Dout[95]), .B(Dout[94]), .Y(
        \U1/aes_core/SB1/n2540 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U612  ( .A(Dout[93]), .B(Dout[92]), .Y(
        \U1/aes_core/SB1/n2531 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U611  ( .A(\U1/aes_core/SB1/n2540 ), .B(
        \U1/aes_core/SB1/n2531 ), .Y(\U1/aes_core/SB1/n2604 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U610  ( .A(Dout[89]), .Y(
        \U1/aes_core/SB1/n2525 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U609  ( .A(Dout[88]), .Y(
        \U1/aes_core/SB1/n2522 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U608  ( .A(\U1/aes_core/SB1/n2525 ), .B(
        \U1/aes_core/SB1/n2522 ), .Y(\U1/aes_core/SB1/n2532 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U607  ( .A(Dout[91]), .B(Dout[90]), .Y(
        \U1/aes_core/SB1/n2552 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U606  ( .A(\U1/aes_core/SB1/n2532 ), .B(
        \U1/aes_core/SB1/n2552 ), .Y(\U1/aes_core/SB1/n2907 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U605  ( .A(\U1/aes_core/SB1/n2604 ), .B(
        \U1/aes_core/SB1/n2907 ), .Y(\U1/aes_core/SB1/n2693 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U604  ( .A(Dout[90]), .B(Dout[91]), .Y(
        \U1/aes_core/SB1/n2535 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U603  ( .A(\U1/aes_core/SB1/n2535 ), .B(
        \U1/aes_core/SB1/n2532 ), .Y(\U1/aes_core/SB1/n2824 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U602  ( .A(Dout[95]), .Y(
        \U1/aes_core/SB1/n2528 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U601  ( .A(\U1/aes_core/SB1/n2528 ), .B(
        Dout[94]), .Y(\U1/aes_core/SB1/n2558 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U600  ( .A(\U1/aes_core/SB1/n2558 ), .B(
        \U1/aes_core/SB1/n2531 ), .Y(\U1/aes_core/SB1/n2603 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U599  ( .A(\U1/aes_core/SB1/n2824 ), .B(
        \U1/aes_core/SB1/n2603 ), .Y(\U1/aes_core/SB1/n2790 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U598  ( .A(Dout[91]), .Y(
        \U1/aes_core/SB1/n2523 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB1/U597  ( .A(Dout[90]), .B(
        \U1/aes_core/SB1/n2523 ), .Y(\U1/aes_core/SB1/n2533 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U596  ( .A(\U1/aes_core/SB1/n2532 ), .B(
        \U1/aes_core/SB1/n2533 ), .Y(\U1/aes_core/SB1/n2755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U595  ( .A(\U1/aes_core/SB1/n2755 ), .Y(
        \U1/aes_core/SB1/n2941 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U594  ( .A(Dout[92]), .Y(
        \U1/aes_core/SB1/n2524 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U593  ( .A(\U1/aes_core/SB1/n2524 ), .B(
        Dout[93]), .Y(\U1/aes_core/SB1/n2539 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U592  ( .A(Dout[94]), .Y(
        \U1/aes_core/SB1/n2527 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U591  ( .A(\U1/aes_core/SB1/n2527 ), .B(
        Dout[95]), .Y(\U1/aes_core/SB1/n2549 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U590  ( .A(\U1/aes_core/SB1/n2539 ), .B(
        \U1/aes_core/SB1/n2549 ), .Y(\U1/aes_core/SB1/n2776 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U589  ( .A(\U1/aes_core/SB1/n2776 ), .Y(
        \U1/aes_core/SB1/n2874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U588  ( .A(\U1/aes_core/SB1/n2941 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2733 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U587  ( .A(\U1/aes_core/SB1/n2604 ), .Y(
        \U1/aes_core/SB1/n2910 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U586  ( .A(Dout[89]), .B(Dout[88]), .Y(
        \U1/aes_core/SB1/n2536 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U585  ( .A(\U1/aes_core/SB1/n2536 ), .B(
        \U1/aes_core/SB1/n2552 ), .Y(\U1/aes_core/SB1/n2842 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U584  ( .A(\U1/aes_core/SB1/n2842 ), .Y(
        \U1/aes_core/SB1/n2951 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U583  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2951 ), .Y(\U1/aes_core/SB1/n2847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U582  ( .A(\U1/aes_core/SB1/n2522 ), .B(
        Dout[89]), .Y(\U1/aes_core/SB1/n2551 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U581  ( .A(\U1/aes_core/SB1/n2533 ), .B(
        \U1/aes_core/SB1/n2551 ), .Y(\U1/aes_core/SB1/n2742 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U580  ( .A(\U1/aes_core/SB1/n2742 ), .Y(
        \U1/aes_core/SB1/n2831 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U579  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2711 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U578  ( .A(\U1/aes_core/SB1/n2733 ), .B(
        \U1/aes_core/SB1/n2847 ), .C(\U1/aes_core/SB1/n2711 ), .Y(
        \U1/aes_core/SB1/n2571 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U577  ( .A(\U1/aes_core/SB1/n2531 ), .B(
        \U1/aes_core/SB1/n2549 ), .Y(\U1/aes_core/SB1/n2775 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U576  ( .A(\U1/aes_core/SB1/n2523 ), .B(
        Dout[90]), .Y(\U1/aes_core/SB1/n2542 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U575  ( .A(\U1/aes_core/SB1/n2542 ), .B(
        \U1/aes_core/SB1/n2551 ), .Y(\U1/aes_core/SB1/n2773 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U574  ( .A(\U1/aes_core/SB1/n2775 ), .B(
        \U1/aes_core/SB1/n2773 ), .Y(\U1/aes_core/SB1/n2688 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U573  ( .A(\U1/aes_core/SB1/n2603 ), .Y(
        \U1/aes_core/SB1/n2912 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U572  ( .A(Dout[93]), .Y(
        \U1/aes_core/SB1/n2526 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U571  ( .A(\U1/aes_core/SB1/n2524 ), .B(
        \U1/aes_core/SB1/n2526 ), .Y(\U1/aes_core/SB1/n2550 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U570  ( .A(\U1/aes_core/SB1/n2540 ), .B(
        \U1/aes_core/SB1/n2550 ), .Y(\U1/aes_core/SB1/n2955 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U569  ( .A(\U1/aes_core/SB1/n2955 ), .Y(
        \U1/aes_core/SB1/n2865 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U568  ( .A(\U1/aes_core/SB1/n2525 ), .B(
        Dout[88]), .Y(\U1/aes_core/SB1/n2541 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U567  ( .A(\U1/aes_core/SB1/n2541 ), .B(
        \U1/aes_core/SB1/n2552 ), .Y(\U1/aes_core/SB1/n2920 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U566  ( .A(\U1/aes_core/SB1/n2920 ), .Y(
        \U1/aes_core/SB1/n2747 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U565  ( .A0(\U1/aes_core/SB1/n2912 ), 
        .A1(\U1/aes_core/SB1/n2865 ), .B0(\U1/aes_core/SB1/n2747 ), .Y(
        \U1/aes_core/SB1/n2530 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U564  ( .A(\U1/aes_core/SB1/n2536 ), .B(
        \U1/aes_core/SB1/n2533 ), .Y(\U1/aes_core/SB1/n2908 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U563  ( .A(\U1/aes_core/SB1/n2908 ), .Y(
        \U1/aes_core/SB1/n2873 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U562  ( .A(\U1/aes_core/SB1/n2526 ), .B(
        Dout[92]), .Y(\U1/aes_core/SB1/n2557 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U561  ( .A(\U1/aes_core/SB1/n2549 ), .B(
        \U1/aes_core/SB1/n2557 ), .Y(\U1/aes_core/SB1/n2948 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U560  ( .A(\U1/aes_core/SB1/n2775 ), .B(
        \U1/aes_core/SB1/n2948 ), .Y(\U1/aes_core/SB1/n2666 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U559  ( .A(\U1/aes_core/SB1/n2528 ), .B(
        \U1/aes_core/SB1/n2527 ), .Y(\U1/aes_core/SB1/n2548 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U558  ( .A(\U1/aes_core/SB1/n2539 ), .B(
        \U1/aes_core/SB1/n2548 ), .Y(\U1/aes_core/SB1/n2923 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U557  ( .A(\U1/aes_core/SB1/n2923 ), .Y(
        \U1/aes_core/SB1/n2647 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U556  ( .A0(\U1/aes_core/SB1/n2873 ), 
        .A1(\U1/aes_core/SB1/n2666 ), .B0(\U1/aes_core/SB1/n2647 ), .B1(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2529 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U555  ( .AN(\U1/aes_core/SB1/n2688 ), 
        .B(\U1/aes_core/SB1/n2530 ), .C(\U1/aes_core/SB1/n2529 ), .Y(
        \U1/aes_core/SB1/n2570 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U554  ( .A(\U1/aes_core/SB1/n2531 ), .B(
        \U1/aes_core/SB1/n2548 ), .Y(\U1/aes_core/SB1/n2792 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U553  ( .A(\U1/aes_core/SB1/n2535 ), .B(
        \U1/aes_core/SB1/n2536 ), .Y(\U1/aes_core/SB1/n2958 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U552  ( .A(\U1/aes_core/SB1/n2558 ), .B(
        \U1/aes_core/SB1/n2539 ), .Y(\U1/aes_core/SB1/n2843 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U551  ( .A(\U1/aes_core/SB1/n2535 ), .B(
        \U1/aes_core/SB1/n2541 ), .Y(\U1/aes_core/SB1/n2840 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U550  ( .A(\U1/aes_core/SB1/n2532 ), .B(
        \U1/aes_core/SB1/n2542 ), .Y(\U1/aes_core/SB1/n2845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U549  ( .A(\U1/aes_core/SB1/n2845 ), .Y(
        \U1/aes_core/SB1/n2825 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U548  ( .A(\U1/aes_core/SB1/n2948 ), .Y(
        \U1/aes_core/SB1/n2661 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U547  ( .A(\U1/aes_core/SB1/n2533 ), .B(
        \U1/aes_core/SB1/n2541 ), .Y(\U1/aes_core/SB1/n2863 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U546  ( .A(\U1/aes_core/SB1/n2863 ), .Y(
        \U1/aes_core/SB1/n2909 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U545  ( .A0(\U1/aes_core/SB1/n2825 ), 
        .A1(\U1/aes_core/SB1/n2910 ), .B0(\U1/aes_core/SB1/n2661 ), .B1(
        \U1/aes_core/SB1/n2909 ), .Y(\U1/aes_core/SB1/n2534 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U544  ( .A0(\U1/aes_core/SB1/n2792 ), 
        .A1(\U1/aes_core/SB1/n2958 ), .B0(\U1/aes_core/SB1/n2843 ), .B1(
        \U1/aes_core/SB1/n2840 ), .C0(\U1/aes_core/SB1/n2534 ), .Y(
        \U1/aes_core/SB1/n2569 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U543  ( .A(\U1/aes_core/SB1/n2845 ), .B(
        \U1/aes_core/SB1/n2792 ), .Y(\U1/aes_core/SB1/n2654 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U542  ( .A(\U1/aes_core/SB1/n2840 ), .B(
        \U1/aes_core/SB1/n2775 ), .Y(\U1/aes_core/SB1/n2664 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U541  ( .A(\U1/aes_core/SB1/n2664 ), .Y(
        \U1/aes_core/SB1/n2538 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U540  ( .A(\U1/aes_core/SB1/n2535 ), .B(
        \U1/aes_core/SB1/n2551 ), .Y(\U1/aes_core/SB1/n2936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U539  ( .A(\U1/aes_core/SB1/n2936 ), .Y(
        \U1/aes_core/SB1/n2864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U538  ( .A(\U1/aes_core/SB1/n2536 ), .B(
        \U1/aes_core/SB1/n2542 ), .Y(\U1/aes_core/SB1/n2921 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U537  ( .A(\U1/aes_core/SB1/n2921 ), .Y(
        \U1/aes_core/SB1/n2932 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U536  ( .A0(\U1/aes_core/SB1/n2864 ), 
        .A1(\U1/aes_core/SB1/n2932 ), .B0(\U1/aes_core/SB1/n2865 ), .Y(
        \U1/aes_core/SB1/n2537 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U535  ( .A(\U1/aes_core/SB1/n2540 ), .B(
        \U1/aes_core/SB1/n2557 ), .Y(\U1/aes_core/SB1/n2937 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U534  ( .A(\U1/aes_core/SB1/n2937 ), .Y(
        \U1/aes_core/SB1/n2866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U533  ( .A(\U1/aes_core/SB1/n2866 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2681 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U532  ( .AN(\U1/aes_core/SB1/n2654 ), 
        .B(\U1/aes_core/SB1/n2538 ), .C(\U1/aes_core/SB1/n2537 ), .D(
        \U1/aes_core/SB1/n2681 ), .Y(\U1/aes_core/SB1/n2547 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U531  ( .A(\U1/aes_core/SB1/n2550 ), .B(
        \U1/aes_core/SB1/n2548 ), .Y(\U1/aes_core/SB1/n2957 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U530  ( .A(\U1/aes_core/SB1/n2540 ), .B(
        \U1/aes_core/SB1/n2539 ), .Y(\U1/aes_core/SB1/n2949 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U529  ( .A0(\U1/aes_core/SB1/n2603 ), 
        .A1(\U1/aes_core/SB1/n2755 ), .B0(\U1/aes_core/SB1/n2957 ), .B1(
        \U1/aes_core/SB1/n2845 ), .C0(\U1/aes_core/SB1/n2949 ), .C1(
        \U1/aes_core/SB1/n2863 ), .Y(\U1/aes_core/SB1/n2546 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U528  ( .A(\U1/aes_core/SB1/n2908 ), .B(
        \U1/aes_core/SB1/n2603 ), .Y(\U1/aes_core/SB1/n2739 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U527  ( .A(\U1/aes_core/SB1/n2661 ), .B(
        \U1/aes_core/SB1/n2825 ), .Y(\U1/aes_core/SB1/n2692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U526  ( .A(\U1/aes_core/SB1/n2909 ), .B(
        \U1/aes_core/SB1/n2910 ), .Y(\U1/aes_core/SB1/n2712 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U525  ( .A(\U1/aes_core/SB1/n2843 ), .Y(
        \U1/aes_core/SB1/n2938 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U524  ( .A(\U1/aes_core/SB1/n2938 ), .B(
        \U1/aes_core/SB1/n2747 ), .Y(\U1/aes_core/SB1/n2750 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U523  ( .AN(\U1/aes_core/SB1/n2739 ), 
        .B(\U1/aes_core/SB1/n2692 ), .C(\U1/aes_core/SB1/n2712 ), .D(
        \U1/aes_core/SB1/n2750 ), .Y(\U1/aes_core/SB1/n2545 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U522  ( .A(\U1/aes_core/SB1/n2558 ), .B(
        \U1/aes_core/SB1/n2550 ), .Y(\U1/aes_core/SB1/n2662 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U521  ( .A(\U1/aes_core/SB1/n2662 ), .B(
        \U1/aes_core/SB1/n2920 ), .Y(\U1/aes_core/SB1/n2816 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U520  ( .A(\U1/aes_core/SB1/n2542 ), .B(
        \U1/aes_core/SB1/n2541 ), .Y(\U1/aes_core/SB1/n2956 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U519  ( .A(\U1/aes_core/SB1/n2923 ), .B(
        \U1/aes_core/SB1/n2956 ), .Y(\U1/aes_core/SB1/n2781 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U518  ( .A(\U1/aes_core/SB1/n2781 ), .Y(
        \U1/aes_core/SB1/n2543 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U517  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2747 ), .Y(\U1/aes_core/SB1/n2800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U516  ( .A(\U1/aes_core/SB1/n2956 ), .Y(
        \U1/aes_core/SB1/n2939 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U515  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2939 ), .Y(\U1/aes_core/SB1/n2851 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U514  ( .AN(\U1/aes_core/SB1/n2816 ), 
        .B(\U1/aes_core/SB1/n2543 ), .C(\U1/aes_core/SB1/n2800 ), .D(
        \U1/aes_core/SB1/n2851 ), .Y(\U1/aes_core/SB1/n2544 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U513  ( .A(\U1/aes_core/SB1/n2547 ), .B(
        \U1/aes_core/SB1/n2546 ), .C(\U1/aes_core/SB1/n2545 ), .D(
        \U1/aes_core/SB1/n2544 ), .Y(\U1/aes_core/SB1/n2643 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U512  ( .A(\U1/aes_core/SB1/n2842 ), .B(
        \U1/aes_core/SB1/n2662 ), .Y(\U1/aes_core/SB1/n2850 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U511  ( .A(\U1/aes_core/SB1/n2557 ), .B(
        \U1/aes_core/SB1/n2548 ), .Y(\U1/aes_core/SB1/n2758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U510  ( .A(\U1/aes_core/SB1/n2824 ), .B(
        \U1/aes_core/SB1/n2758 ), .Y(\U1/aes_core/SB1/n2729 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U509  ( .A(\U1/aes_core/SB1/n2957 ), .Y(
        \U1/aes_core/SB1/n2913 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U508  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2873 ), .Y(\U1/aes_core/SB1/n2678 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U507  ( .A0(\U1/aes_core/SB1/n2758 ), 
        .A1(\U1/aes_core/SB1/n2956 ), .B0(\U1/aes_core/SB1/n2678 ), .Y(
        \U1/aes_core/SB1/n2556 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U506  ( .A(\U1/aes_core/SB1/n2773 ), .Y(
        \U1/aes_core/SB1/n2868 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U505  ( .A(\U1/aes_core/SB1/n2868 ), .B(
        \U1/aes_core/SB1/n2912 ), .Y(\U1/aes_core/SB1/n2869 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U504  ( .A(\U1/aes_core/SB1/n2912 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2828 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U503  ( .A(\U1/aes_core/SB1/n2550 ), .B(
        \U1/aes_core/SB1/n2549 ), .Y(\U1/aes_core/SB1/n2919 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U502  ( .A(\U1/aes_core/SB1/n2919 ), .Y(
        \U1/aes_core/SB1/n2673 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U501  ( .A(\U1/aes_core/SB1/n2864 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2697 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U500  ( .A(\U1/aes_core/SB1/n2907 ), .Y(
        \U1/aes_core/SB1/n2867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U499  ( .A(\U1/aes_core/SB1/n2867 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2761 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U498  ( .A(\U1/aes_core/SB1/n2869 ), .B(
        \U1/aes_core/SB1/n2828 ), .C(\U1/aes_core/SB1/n2697 ), .D(
        \U1/aes_core/SB1/n2761 ), .Y(\U1/aes_core/SB1/n2555 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U497  ( .A(\U1/aes_core/SB1/n2909 ), .B(
        \U1/aes_core/SB1/n2866 ), .Y(\U1/aes_core/SB1/n2795 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U496  ( .A(\U1/aes_core/SB1/n2951 ), .B(
        \U1/aes_core/SB1/n2866 ), .Y(\U1/aes_core/SB1/n2786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U495  ( .A(\U1/aes_core/SB1/n2949 ), .Y(
        \U1/aes_core/SB1/n2942 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U494  ( .A(\U1/aes_core/SB1/n2825 ), .B(
        \U1/aes_core/SB1/n2942 ), .Y(\U1/aes_core/SB1/n2658 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U493  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2864 ), .Y(\U1/aes_core/SB1/n2769 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U492  ( .A(\U1/aes_core/SB1/n2795 ), .B(
        \U1/aes_core/SB1/n2786 ), .C(\U1/aes_core/SB1/n2658 ), .D(
        \U1/aes_core/SB1/n2769 ), .Y(\U1/aes_core/SB1/n2554 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U491  ( .A(\U1/aes_core/SB1/n2840 ), .Y(
        \U1/aes_core/SB1/n2809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U490  ( .A(\U1/aes_core/SB1/n2661 ), .B(
        \U1/aes_core/SB1/n2809 ), .Y(\U1/aes_core/SB1/n2645 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U489  ( .A(\U1/aes_core/SB1/n2552 ), .B(
        \U1/aes_core/SB1/n2551 ), .Y(\U1/aes_core/SB1/n2875 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U488  ( .A(\U1/aes_core/SB1/n2875 ), .Y(
        \U1/aes_core/SB1/n2930 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U487  ( .A(\U1/aes_core/SB1/n2661 ), .B(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2709 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U486  ( .A(\U1/aes_core/SB1/n2824 ), .Y(
        \U1/aes_core/SB1/n2953 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U485  ( .A(\U1/aes_core/SB1/n2953 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2744 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U484  ( .A(\U1/aes_core/SB1/n2865 ), .B(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2914 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U483  ( .A(\U1/aes_core/SB1/n2645 ), .B(
        \U1/aes_core/SB1/n2709 ), .C(\U1/aes_core/SB1/n2744 ), .D(
        \U1/aes_core/SB1/n2914 ), .Y(\U1/aes_core/SB1/n2553 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U482  ( .A(\U1/aes_core/SB1/n2850 ), .B(
        \U1/aes_core/SB1/n2729 ), .C(\U1/aes_core/SB1/n2556 ), .D(
        \U1/aes_core/SB1/n2555 ), .E(\U1/aes_core/SB1/n2554 ), .F(
        \U1/aes_core/SB1/n2553 ), .Y(\U1/aes_core/SB1/n2632 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U481  ( .A(\U1/aes_core/SB1/n2632 ), .Y(
        \U1/aes_core/SB1/n2567 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U480  ( .A(\U1/aes_core/SB1/n2921 ), .B(
        \U1/aes_core/SB1/n2758 ), .Y(\U1/aes_core/SB1/n2655 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U479  ( .A(\U1/aes_core/SB1/n2558 ), .B(
        \U1/aes_core/SB1/n2557 ), .Y(\U1/aes_core/SB1/n2918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U478  ( .A(\U1/aes_core/SB1/n2918 ), .B(
        \U1/aes_core/SB1/n2773 ), .Y(\U1/aes_core/SB1/n2782 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U477  ( .A(\U1/aes_core/SB1/n2782 ), .Y(
        \U1/aes_core/SB1/n2560 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U476  ( .A(\U1/aes_core/SB1/n2775 ), .Y(
        \U1/aes_core/SB1/n2943 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U475  ( .A0(\U1/aes_core/SB1/n2673 ), 
        .A1(\U1/aes_core/SB1/n2943 ), .B0(\U1/aes_core/SB1/n2930 ), .Y(
        \U1/aes_core/SB1/n2559 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U474  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2809 ), .Y(\U1/aes_core/SB1/n2680 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U473  ( .AN(\U1/aes_core/SB1/n2655 ), 
        .B(\U1/aes_core/SB1/n2560 ), .C(\U1/aes_core/SB1/n2559 ), .D(
        \U1/aes_core/SB1/n2680 ), .Y(\U1/aes_core/SB1/n2564 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U472  ( .A0(\U1/aes_core/SB1/n2907 ), 
        .A1(\U1/aes_core/SB1/n2955 ), .B0(\U1/aes_core/SB1/n2792 ), .B1(
        \U1/aes_core/SB1/n2840 ), .C0(\U1/aes_core/SB1/n2920 ), .C1(
        \U1/aes_core/SB1/n2937 ), .Y(\U1/aes_core/SB1/n2563 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U471  ( .A(\U1/aes_core/SB1/n2955 ), .B(
        \U1/aes_core/SB1/n2958 ), .Y(\U1/aes_core/SB1/n2720 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U470  ( .A(\U1/aes_core/SB1/n2943 ), .B(
        \U1/aes_core/SB1/n2864 ), .Y(\U1/aes_core/SB1/n2853 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U469  ( .A(\U1/aes_core/SB1/n2825 ), .B(
        \U1/aes_core/SB1/n2943 ), .Y(\U1/aes_core/SB1/n2787 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U468  ( .A(\U1/aes_core/SB1/n2809 ), .B(
        \U1/aes_core/SB1/n2910 ), .Y(\U1/aes_core/SB1/n2659 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U467  ( .AN(\U1/aes_core/SB1/n2720 ), 
        .B(\U1/aes_core/SB1/n2853 ), .C(\U1/aes_core/SB1/n2787 ), .D(
        \U1/aes_core/SB1/n2659 ), .Y(\U1/aes_core/SB1/n2562 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U466  ( .A(\U1/aes_core/SB1/n2953 ), .B(
        \U1/aes_core/SB1/n2938 ), .Y(\U1/aes_core/SB1/n2732 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U465  ( .A(\U1/aes_core/SB1/n2809 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U464  ( .A(\U1/aes_core/SB1/n2661 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U463  ( .A(\U1/aes_core/SB1/n2868 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2745 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U462  ( .A(\U1/aes_core/SB1/n2732 ), .B(
        \U1/aes_core/SB1/n2799 ), .C(\U1/aes_core/SB1/n2700 ), .D(
        \U1/aes_core/SB1/n2745 ), .Y(\U1/aes_core/SB1/n2561 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U461  ( .A(\U1/aes_core/SB1/n2564 ), .B(
        \U1/aes_core/SB1/n2563 ), .C(\U1/aes_core/SB1/n2562 ), .D(
        \U1/aes_core/SB1/n2561 ), .Y(\U1/aes_core/SB1/n2565 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U460  ( .A(\U1/aes_core/SB1/n2565 ), .Y(
        \U1/aes_core/SB1/n2935 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U459  ( .A(\U1/aes_core/SB1/n2951 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2566 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U458  ( .AN(\U1/aes_core/SB1/n2643 ), 
        .B(\U1/aes_core/SB1/n2567 ), .C(\U1/aes_core/SB1/n2935 ), .D(
        \U1/aes_core/SB1/n2566 ), .Y(\U1/aes_core/SB1/n2568 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U457  ( .A(\U1/aes_core/SB1/n2693 ), .B(
        \U1/aes_core/SB1/n2790 ), .C(\U1/aes_core/SB1/n2571 ), .D(
        \U1/aes_core/SB1/n2570 ), .E(\U1/aes_core/SB1/n2569 ), .F(
        \U1/aes_core/SB1/n2568 ), .Y(\U1/aes_core/SB1/n2622 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U456  ( .A(\U1/aes_core/SB1/n2936 ), .B(
        \U1/aes_core/SB1/n2603 ), .Y(\U1/aes_core/SB1/n2738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U455  ( .A(\U1/aes_core/SB1/n2865 ), .B(
        \U1/aes_core/SB1/n2953 ), .Y(\U1/aes_core/SB1/n2789 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U454  ( .A(\U1/aes_core/SB1/n2942 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2691 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U453  ( .A(\U1/aes_core/SB1/n2662 ), .Y(
        \U1/aes_core/SB1/n2931 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U452  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2714 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U451  ( .AN(\U1/aes_core/SB1/n2738 ), 
        .B(\U1/aes_core/SB1/n2789 ), .C(\U1/aes_core/SB1/n2691 ), .D(
        \U1/aes_core/SB1/n2714 ), .Y(\U1/aes_core/SB1/n2578 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U450  ( .A(\U1/aes_core/SB1/n2923 ), .B(
        \U1/aes_core/SB1/n2773 ), .Y(\U1/aes_core/SB1/n2815 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U449  ( .A(\U1/aes_core/SB1/n2825 ), .B(
        \U1/aes_core/SB1/n2912 ), .Y(\U1/aes_core/SB1/n2671 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U448  ( .A0(\U1/aes_core/SB1/n2932 ), 
        .A1(\U1/aes_core/SB1/n2831 ), .B0(\U1/aes_core/SB1/n2661 ), .Y(
        \U1/aes_core/SB1/n2572 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U447  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2763 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U446  ( .AN(\U1/aes_core/SB1/n2815 ), 
        .B(\U1/aes_core/SB1/n2671 ), .C(\U1/aes_core/SB1/n2572 ), .D(
        \U1/aes_core/SB1/n2763 ), .Y(\U1/aes_core/SB1/n2573 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U445  ( .A(\U1/aes_core/SB1/n2573 ), .Y(
        \U1/aes_core/SB1/n2577 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U444  ( .A(\U1/aes_core/SB1/n2792 ), .Y(
        \U1/aes_core/SB1/n2933 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U443  ( .A(\U1/aes_core/SB1/n2958 ), .Y(
        \U1/aes_core/SB1/n2832 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U442  ( .A0(\U1/aes_core/SB1/n2953 ), 
        .A1(\U1/aes_core/SB1/n2866 ), .B0(\U1/aes_core/SB1/n2933 ), .B1(
        \U1/aes_core/SB1/n2747 ), .C0(\U1/aes_core/SB1/n2832 ), .C1(
        \U1/aes_core/SB1/n2931 ), .Y(\U1/aes_core/SB1/n2576 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U441  ( .A0(\U1/aes_core/SB1/n2758 ), 
        .A1(\U1/aes_core/SB1/n2936 ), .B0(\U1/aes_core/SB1/n2956 ), .B1(
        \U1/aes_core/SB1/n2957 ), .Y(\U1/aes_core/SB1/n2574 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U440  ( .A0(\U1/aes_core/SB1/n2809 ), 
        .A1(\U1/aes_core/SB1/n2647 ), .B0(\U1/aes_core/SB1/n2865 ), .B1(
        \U1/aes_core/SB1/n2909 ), .C0(\U1/aes_core/SB1/n2574 ), .Y(
        \U1/aes_core/SB1/n2575 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U439  ( .AN(\U1/aes_core/SB1/n2578 ), 
        .B(\U1/aes_core/SB1/n2577 ), .C(\U1/aes_core/SB1/n2576 ), .D(
        \U1/aes_core/SB1/n2575 ), .Y(\U1/aes_core/SB1/n2641 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U438  ( .A(\U1/aes_core/SB1/n2957 ), .B(
        \U1/aes_core/SB1/n2773 ), .Y(\U1/aes_core/SB1/n2656 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U437  ( .A0(\U1/aes_core/SB1/n2843 ), 
        .A1(\U1/aes_core/SB1/n2957 ), .B0(\U1/aes_core/SB1/n2875 ), .Y(
        \U1/aes_core/SB1/n2583 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U436  ( .A(\U1/aes_core/SB1/n2875 ), .B(
        \U1/aes_core/SB1/n2863 ), .Y(\U1/aes_core/SB1/n2740 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB1/U435  ( .A0(\U1/aes_core/SB1/n2864 ), .A1(
        \U1/aes_core/SB1/n2647 ), .B0(\U1/aes_core/SB1/n2740 ), .B1(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2582 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U434  ( .A0(\U1/aes_core/SB1/n2918 ), 
        .A1(\U1/aes_core/SB1/n2958 ), .B0(\U1/aes_core/SB1/n2662 ), .B1(
        \U1/aes_core/SB1/n2755 ), .C0(\U1/aes_core/SB1/n2920 ), .C1(
        \U1/aes_core/SB1/n2949 ), .Y(\U1/aes_core/SB1/n2581 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U433  ( .A(\U1/aes_core/SB1/n2758 ), .Y(
        \U1/aes_core/SB1/n2826 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U432  ( .A(\U1/aes_core/SB1/n2951 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2852 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U431  ( .A(\U1/aes_core/SB1/n2825 ), .B(
        \U1/aes_core/SB1/n2647 ), .Y(\U1/aes_core/SB1/n2679 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U430  ( .A(\U1/aes_core/SB1/n2661 ), .B(
        \U1/aes_core/SB1/n2868 ), .Y(\U1/aes_core/SB1/n2699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U429  ( .A(\U1/aes_core/SB1/n2825 ), .B(
        \U1/aes_core/SB1/n2866 ), .Y(\U1/aes_core/SB1/n2798 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U428  ( .A(\U1/aes_core/SB1/n2852 ), .B(
        \U1/aes_core/SB1/n2679 ), .C(\U1/aes_core/SB1/n2699 ), .D(
        \U1/aes_core/SB1/n2798 ), .Y(\U1/aes_core/SB1/n2580 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U427  ( .A(\U1/aes_core/SB1/n2845 ), .B(
        \U1/aes_core/SB1/n2758 ), .Y(\U1/aes_core/SB1/n2721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U426  ( .A(\U1/aes_core/SB1/n2831 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2731 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U425  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2747 ), .Y(\U1/aes_core/SB1/n2762 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB1/U424  ( .AN(\U1/aes_core/SB1/n2721 ), 
        .B(\U1/aes_core/SB1/n2731 ), .C(\U1/aes_core/SB1/n2762 ), .Y(
        \U1/aes_core/SB1/n2579 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U423  ( .A(\U1/aes_core/SB1/n2656 ), .B(
        \U1/aes_core/SB1/n2583 ), .C(\U1/aes_core/SB1/n2582 ), .D(
        \U1/aes_core/SB1/n2581 ), .E(\U1/aes_core/SB1/n2580 ), .F(
        \U1/aes_core/SB1/n2579 ), .Y(\U1/aes_core/SB1/n2964 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U422  ( .A0(\U1/aes_core/SB1/n2661 ), 
        .A1(\U1/aes_core/SB1/n2910 ), .B0(\U1/aes_core/SB1/n2941 ), .Y(
        \U1/aes_core/SB1/n2584 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U421  ( .A(\U1/aes_core/SB1/n2647 ), .B(
        \U1/aes_core/SB1/n2747 ), .Y(\U1/aes_core/SB1/n2784 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U420  ( .A(\U1/aes_core/SB1/n2864 ), .B(
        \U1/aes_core/SB1/n2933 ), .Y(\U1/aes_core/SB1/n2676 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U419  ( .A(\U1/aes_core/SB1/n2933 ), .B(
        \U1/aes_core/SB1/n2868 ), .Y(\U1/aes_core/SB1/n2727 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U418  ( .A(\U1/aes_core/SB1/n2584 ), .B(
        \U1/aes_core/SB1/n2784 ), .C(\U1/aes_core/SB1/n2676 ), .D(
        \U1/aes_core/SB1/n2727 ), .Y(\U1/aes_core/SB1/n2588 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U417  ( .A0(\U1/aes_core/SB1/n2936 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2662 ), .B1(
        \U1/aes_core/SB1/n2908 ), .C0(\U1/aes_core/SB1/n2937 ), .C1(
        \U1/aes_core/SB1/n2773 ), .Y(\U1/aes_core/SB1/n2587 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U416  ( .A(\U1/aes_core/SB1/n2867 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U415  ( .A(\U1/aes_core/SB1/n2866 ), .B(
        \U1/aes_core/SB1/n2939 ), .Y(\U1/aes_core/SB1/n2848 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U414  ( .A(\U1/aes_core/SB1/n2866 ), .B(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2695 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U413  ( .A(\U1/aes_core/SB1/n2942 ), .B(
        \U1/aes_core/SB1/n2932 ), .Y(\U1/aes_core/SB1/n2657 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U412  ( .A(\U1/aes_core/SB1/n2708 ), .B(
        \U1/aes_core/SB1/n2848 ), .C(\U1/aes_core/SB1/n2695 ), .D(
        \U1/aes_core/SB1/n2657 ), .Y(\U1/aes_core/SB1/n2586 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U411  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2770 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U410  ( .A(\U1/aes_core/SB1/n2951 ), .B(
        \U1/aes_core/SB1/n2912 ), .Y(\U1/aes_core/SB1/n2743 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U409  ( .A(\U1/aes_core/SB1/n2941 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2794 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U408  ( .A(\U1/aes_core/SB1/n2673 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2644 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U407  ( .A(\U1/aes_core/SB1/n2770 ), .B(
        \U1/aes_core/SB1/n2743 ), .C(\U1/aes_core/SB1/n2794 ), .D(
        \U1/aes_core/SB1/n2644 ), .Y(\U1/aes_core/SB1/n2585 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U406  ( .A(\U1/aes_core/SB1/n2588 ), .B(
        \U1/aes_core/SB1/n2587 ), .C(\U1/aes_core/SB1/n2586 ), .D(
        \U1/aes_core/SB1/n2585 ), .Y(\U1/aes_core/SB1/n2630 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U405  ( .A(\U1/aes_core/SB1/n2622 ), .B(
        \U1/aes_core/SB1/n2641 ), .C(\U1/aes_core/SB1/n2964 ), .D(
        \U1/aes_core/SB1/n2630 ), .Y(\U1/aes_core/SB1/n2597 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U404  ( .A(\U1/aes_core/SB1/n2918 ), .Y(
        \U1/aes_core/SB1/n2821 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U403  ( .A0(\U1/aes_core/SB1/n2773 ), 
        .A1(\U1/aes_core/SB1/n2604 ), .B0(\U1/aes_core/SB1/n2742 ), .B1(
        \U1/aes_core/SB1/n2949 ), .Y(\U1/aes_core/SB1/n2589 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U402  ( .A0(\U1/aes_core/SB1/n2821 ), 
        .A1(\U1/aes_core/SB1/n2873 ), .B0(\U1/aes_core/SB1/n2943 ), .B1(
        \U1/aes_core/SB1/n2951 ), .C0(\U1/aes_core/SB1/n2589 ), .Y(
        \U1/aes_core/SB1/n2596 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U401  ( .A(\U1/aes_core/SB1/n2842 ), .B(
        \U1/aes_core/SB1/n2845 ), .Y(\U1/aes_core/SB1/n2841 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U400  ( .A0(\U1/aes_core/SB1/n2776 ), 
        .A1(\U1/aes_core/SB1/n2845 ), .B0(\U1/aes_core/SB1/n2758 ), .B1(
        \U1/aes_core/SB1/n2907 ), .Y(\U1/aes_core/SB1/n2590 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U399  ( .A0(\U1/aes_core/SB1/n2673 ), 
        .A1(\U1/aes_core/SB1/n2841 ), .B0(\U1/aes_core/SB1/n2913 ), .B1(
        \U1/aes_core/SB1/n2932 ), .C0(\U1/aes_core/SB1/n2590 ), .Y(
        \U1/aes_core/SB1/n2595 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U398  ( .A(\U1/aes_core/SB1/n2937 ), .B(
        \U1/aes_core/SB1/n2775 ), .Y(\U1/aes_core/SB1/n2593 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U397  ( .A(\U1/aes_core/SB1/n2866 ), .B(
        \U1/aes_core/SB1/n2912 ), .Y(\U1/aes_core/SB1/n2833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U396  ( .A(\U1/aes_core/SB1/n2833 ), .Y(
        \U1/aes_core/SB1/n2592 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U395  ( .A(\U1/aes_core/SB1/n2824 ), .B(
        \U1/aes_core/SB1/n2918 ), .Y(\U1/aes_core/SB1/n2705 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U394  ( .A(\U1/aes_core/SB1/n2923 ), .B(
        \U1/aes_core/SB1/n2921 ), .Y(\U1/aes_core/SB1/n2858 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U392  ( .A(\U1/aes_core/SB1/n2873 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2715 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U390  ( .A0(\U1/aes_core/SB1/n2832 ), 
        .A1(\U1/aes_core/SB1/n2593 ), .B0(\U1/aes_core/SB1/n2809 ), .B1(
        \U1/aes_core/SB1/n2592 ), .C0(\U1/aes_core/SB1/n2591 ), .Y(
        \U1/aes_core/SB1/n2594 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U389  ( .AN(\U1/aes_core/SB1/n2597 ), 
        .B(\U1/aes_core/SB1/n2596 ), .C(\U1/aes_core/SB1/n2595 ), .D(
        \U1/aes_core/SB1/n2594 ), .Y(\U1/aes_core/sb1 [24]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U388  ( .A(\U1/aes_core/SB1/n2845 ), .B(
        \U1/aes_core/SB1/n2662 ), .Y(\U1/aes_core/SB1/n2722 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U387  ( .A(\U1/aes_core/SB1/n2792 ), .B(
        \U1/aes_core/SB1/n2842 ), .Y(\U1/aes_core/SB1/n2682 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U386  ( .A(\U1/aes_core/SB1/n2809 ), .B(
        \U1/aes_core/SB1/n2941 ), .Y(\U1/aes_core/SB1/n2791 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U385  ( .A0(\U1/aes_core/SB1/n2791 ), 
        .A1(\U1/aes_core/SB1/n2845 ), .B0(\U1/aes_core/SB1/n2955 ), .Y(
        \U1/aes_core/SB1/n2602 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U384  ( .A(\U1/aes_core/SB1/n2873 ), .B(
        \U1/aes_core/SB1/n2942 ), .Y(\U1/aes_core/SB1/n2698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U383  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2873 ), .Y(\U1/aes_core/SB1/n2797 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U382  ( .A(\U1/aes_core/SB1/n2939 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2730 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U381  ( .A(\U1/aes_core/SB1/n2698 ), .B(
        \U1/aes_core/SB1/n2797 ), .C(\U1/aes_core/SB1/n2730 ), .Y(
        \U1/aes_core/SB1/n2601 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U380  ( .A(\U1/aes_core/SB1/n2873 ), .B(
        \U1/aes_core/SB1/n2953 ), .Y(\U1/aes_core/SB1/n2757 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U379  ( .A(\U1/aes_core/SB1/n2939 ), .B(
        \U1/aes_core/SB1/n2930 ), .C(\U1/aes_core/SB1/n2951 ), .Y(
        \U1/aes_core/SB1/n2598 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U378  ( .A0(\U1/aes_core/SB1/n2757 ), 
        .A1(\U1/aes_core/SB1/n2919 ), .B0(\U1/aes_core/SB1/n2598 ), .B1(
        \U1/aes_core/SB1/n2949 ), .C0(\U1/aes_core/SB1/n2792 ), .C1(
        \U1/aes_core/SB1/n2824 ), .Y(\U1/aes_core/SB1/n2600 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U377  ( .A0(\U1/aes_core/SB1/n2920 ), 
        .A1(\U1/aes_core/SB1/n2948 ), .B0(\U1/aes_core/SB1/n2921 ), .B1(
        \U1/aes_core/SB1/n2918 ), .Y(\U1/aes_core/SB1/n2599 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U376  ( .A(\U1/aes_core/SB1/n2722 ), .B(
        \U1/aes_core/SB1/n2682 ), .C(\U1/aes_core/SB1/n2602 ), .D(
        \U1/aes_core/SB1/n2601 ), .E(\U1/aes_core/SB1/n2600 ), .F(
        \U1/aes_core/SB1/n2599 ), .Y(\U1/aes_core/SB1/n2963 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U375  ( .A(\U1/aes_core/SB1/n2773 ), .B(
        \U1/aes_core/SB1/n2758 ), .Y(\U1/aes_core/SB1/n2648 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U374  ( .A0(\U1/aes_core/SB1/n2773 ), 
        .A1(\U1/aes_core/SB1/n2863 ), .B0(\U1/aes_core/SB1/n2662 ), .Y(
        \U1/aes_core/SB1/n2609 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U373  ( .A(\U1/aes_core/SB1/n2867 ), .B(
        \U1/aes_core/SB1/n2873 ), .Y(\U1/aes_core/SB1/n2650 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U372  ( .A0(\U1/aes_core/SB1/n2755 ), 
        .A1(\U1/aes_core/SB1/n2923 ), .B0(\U1/aes_core/SB1/n2650 ), .B1(
        \U1/aes_core/SB1/n2937 ), .Y(\U1/aes_core/SB1/n2608 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U371  ( .A0(\U1/aes_core/SB1/n2742 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2907 ), .B1(
        \U1/aes_core/SB1/n2792 ), .C0(\U1/aes_core/SB1/n2921 ), .C1(
        \U1/aes_core/SB1/n2843 ), .Y(\U1/aes_core/SB1/n2607 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U370  ( .A(\U1/aes_core/SB1/n2956 ), .B(
        \U1/aes_core/SB1/n2603 ), .Y(\U1/aes_core/SB1/n2706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U369  ( .A(\U1/aes_core/SB1/n2943 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U368  ( .A(\U1/aes_core/SB1/n2864 ), .B(
        \U1/aes_core/SB1/n2938 ), .Y(\U1/aes_core/SB1/n2723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U367  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2953 ), .Y(\U1/aes_core/SB1/n2827 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U366  ( .AN(\U1/aes_core/SB1/n2706 ), 
        .B(\U1/aes_core/SB1/n2713 ), .C(\U1/aes_core/SB1/n2723 ), .D(
        \U1/aes_core/SB1/n2827 ), .Y(\U1/aes_core/SB1/n2606 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U365  ( .A(\U1/aes_core/SB1/n2824 ), .B(
        \U1/aes_core/SB1/n2604 ), .Y(\U1/aes_core/SB1/n2806 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U364  ( .A(\U1/aes_core/SB1/n2923 ), .B(
        \U1/aes_core/SB1/n2907 ), .Y(\U1/aes_core/SB1/n2859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U362  ( .A(\U1/aes_core/SB1/n2647 ), .B(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2672 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U360  ( .A(\U1/aes_core/SB1/n2648 ), .B(
        \U1/aes_core/SB1/n2609 ), .C(\U1/aes_core/SB1/n2608 ), .D(
        \U1/aes_core/SB1/n2607 ), .E(\U1/aes_core/SB1/n2606 ), .F(
        \U1/aes_core/SB1/n2605 ), .Y(\U1/aes_core/SB1/n2642 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U359  ( .A(\U1/aes_core/SB1/n2840 ), .B(
        \U1/aes_core/SB1/n2662 ), .Y(\U1/aes_core/SB1/n2660 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U358  ( .A(\U1/aes_core/SB1/n2792 ), .B(
        \U1/aes_core/SB1/n2742 ), .Y(\U1/aes_core/SB1/n2872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U357  ( .A(\U1/aes_core/SB1/n2773 ), .B(
        \U1/aes_core/SB1/n2843 ), .Y(\U1/aes_core/SB1/n2710 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U356  ( .A(\U1/aes_core/SB1/n2958 ), .B(
        \U1/aes_core/SB1/n2843 ), .Y(\U1/aes_core/SB1/n2725 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U355  ( .A(\U1/aes_core/SB1/n2868 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2785 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U354  ( .A(\U1/aes_core/SB1/n2939 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2677 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U353  ( .A(\U1/aes_core/SB1/n2943 ), .B(
        \U1/aes_core/SB1/n2939 ), .Y(\U1/aes_core/SB1/n2771 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U352  ( .A(\U1/aes_core/SB1/n2832 ), .B(
        \U1/aes_core/SB1/n2910 ), .Y(\U1/aes_core/SB1/n2696 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U351  ( .A(\U1/aes_core/SB1/n2785 ), .B(
        \U1/aes_core/SB1/n2677 ), .C(\U1/aes_core/SB1/n2771 ), .D(
        \U1/aes_core/SB1/n2696 ), .Y(\U1/aes_core/SB1/n2613 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U350  ( .A(\U1/aes_core/SB1/n2958 ), .B(
        \U1/aes_core/SB1/n2758 ), .Y(\U1/aes_core/SB1/n2746 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U349  ( .A(\U1/aes_core/SB1/n2957 ), .B(
        \U1/aes_core/SB1/n2742 ), .Y(\U1/aes_core/SB1/n2846 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U348  ( .A(\U1/aes_core/SB1/n2863 ), .B(
        \U1/aes_core/SB1/n2923 ), .Y(\U1/aes_core/SB1/n2796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U347  ( .A(\U1/aes_core/SB1/n2824 ), .B(
        \U1/aes_core/SB1/n2923 ), .Y(\U1/aes_core/SB1/n2646 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U346  ( .A0(\U1/aes_core/SB1/n2923 ), 
        .A1(\U1/aes_core/SB1/n2958 ), .B0(\U1/aes_core/SB1/n2758 ), .B1(
        \U1/aes_core/SB1/n2863 ), .Y(\U1/aes_core/SB1/n2611 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U345  ( .A0(\U1/aes_core/SB1/n2742 ), 
        .A1(\U1/aes_core/SB1/n2955 ), .B0(\U1/aes_core/SB1/n2755 ), .B1(
        \U1/aes_core/SB1/n2792 ), .Y(\U1/aes_core/SB1/n2610 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U344  ( .A(\U1/aes_core/SB1/n2746 ), .B(
        \U1/aes_core/SB1/n2846 ), .C(\U1/aes_core/SB1/n2796 ), .D(
        \U1/aes_core/SB1/n2646 ), .E(\U1/aes_core/SB1/n2611 ), .F(
        \U1/aes_core/SB1/n2610 ), .Y(\U1/aes_core/SB1/n2612 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U343  ( .A(\U1/aes_core/SB1/n2660 ), .B(
        \U1/aes_core/SB1/n2872 ), .C(\U1/aes_core/SB1/n2710 ), .D(
        \U1/aes_core/SB1/n2725 ), .E(\U1/aes_core/SB1/n2613 ), .F(
        \U1/aes_core/SB1/n2612 ), .Y(\U1/aes_core/SB1/n2631 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U342  ( .A0(\U1/aes_core/SB1/n2868 ), 
        .A1(\U1/aes_core/SB1/n2865 ), .B0(\U1/aes_core/SB1/n2942 ), .B1(
        \U1/aes_core/SB1/n2809 ), .C0(\U1/aes_core/SB1/n2631 ), .Y(
        \U1/aes_core/SB1/n2614 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U341  ( .A(\U1/aes_core/SB1/n2614 ), .Y(
        \U1/aes_core/SB1/n2621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U340  ( .A(\U1/aes_core/SB1/n2921 ), .B(
        \U1/aes_core/SB1/n2863 ), .Y(\U1/aes_core/SB1/n2911 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U339  ( .A0(\U1/aes_core/SB1/n2867 ), 
        .A1(\U1/aes_core/SB1/n2911 ), .B0(\U1/aes_core/SB1/n2943 ), .Y(
        \U1/aes_core/SB1/n2617 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U338  ( .A0(\U1/aes_core/SB1/n2832 ), 
        .A1(\U1/aes_core/SB1/n2932 ), .B0(\U1/aes_core/SB1/n2874 ), .Y(
        \U1/aes_core/SB1/n2616 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U337  ( .A0(\U1/aes_core/SB1/n2831 ), 
        .A1(\U1/aes_core/SB1/n2873 ), .B0(\U1/aes_core/SB1/n2938 ), .Y(
        \U1/aes_core/SB1/n2615 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U336  ( .A(\U1/aes_core/SB1/n2864 ), .B(
        \U1/aes_core/SB1/n2931 ), .Y(\U1/aes_core/SB1/n2689 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U335  ( .A(\U1/aes_core/SB1/n2617 ), .B(
        \U1/aes_core/SB1/n2616 ), .C(\U1/aes_core/SB1/n2615 ), .D(
        \U1/aes_core/SB1/n2689 ), .Y(\U1/aes_core/SB1/n2620 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U334  ( .A(\U1/aes_core/SB1/n2930 ), .B(
        \U1/aes_core/SB1/n2825 ), .Y(\U1/aes_core/SB1/n2879 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB1/U333  ( .A(\U1/aes_core/SB1/n2879 ), .B(
        \U1/aes_core/SB1/n2920 ), .C(\U1/aes_core/SB1/n2907 ), .Y(
        \U1/aes_core/SB1/n2618 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U332  ( .A0(\U1/aes_core/SB1/n2863 ), 
        .A1(\U1/aes_core/SB1/n2957 ), .B0(\U1/aes_core/SB1/n2618 ), .B1(
        \U1/aes_core/SB1/n2918 ), .C0(\U1/aes_core/SB1/n2956 ), .C1(
        \U1/aes_core/SB1/n2948 ), .Y(\U1/aes_core/SB1/n2619 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U331  ( .A(\U1/aes_core/SB1/n2963 ), .B(
        \U1/aes_core/SB1/n2642 ), .C(\U1/aes_core/SB1/n2622 ), .D(
        \U1/aes_core/SB1/n2621 ), .E(\U1/aes_core/SB1/n2620 ), .F(
        \U1/aes_core/SB1/n2619 ), .Y(\U1/aes_core/sb1 [25]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U330  ( .A0(\U1/aes_core/SB1/n2912 ), 
        .A1(\U1/aes_core/SB1/n2932 ), .B0(\U1/aes_core/SB1/n2953 ), .B1(
        \U1/aes_core/SB1/n2943 ), .Y(\U1/aes_core/SB1/n2623 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U329  ( .A0(\U1/aes_core/SB1/n2842 ), 
        .A1(\U1/aes_core/SB1/n2957 ), .B0(\U1/aes_core/SB1/n2792 ), .B1(
        \U1/aes_core/SB1/n2863 ), .C0(\U1/aes_core/SB1/n2623 ), .Y(
        \U1/aes_core/SB1/n2629 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U328  ( .A(\U1/aes_core/SB1/n2938 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2726 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U327  ( .A(\U1/aes_core/SB1/n2912 ), .B(
        \U1/aes_core/SB1/n2867 ), .Y(\U1/aes_core/SB1/n2707 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U326  ( .A(\U1/aes_core/SB1/n2932 ), .B(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2675 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U325  ( .A(\U1/aes_core/SB1/n2831 ), .B(
        \U1/aes_core/SB1/n2874 ), .Y(\U1/aes_core/SB1/n2694 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U324  ( .A(\U1/aes_core/SB1/n2726 ), .B(
        \U1/aes_core/SB1/n2707 ), .C(\U1/aes_core/SB1/n2675 ), .D(
        \U1/aes_core/SB1/n2694 ), .Y(\U1/aes_core/SB1/n2628 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U323  ( .A(\U1/aes_core/SB1/n2958 ), .B(
        \U1/aes_core/SB1/n2936 ), .Y(\U1/aes_core/SB1/n2820 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U322  ( .A0(\U1/aes_core/SB1/n2868 ), 
        .A1(\U1/aes_core/SB1/n2820 ), .B0(\U1/aes_core/SB1/n2942 ), .Y(
        \U1/aes_core/SB1/n2626 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U321  ( .A0(\U1/aes_core/SB1/n2939 ), 
        .A1(\U1/aes_core/SB1/n2809 ), .B0(\U1/aes_core/SB1/n2821 ), .Y(
        \U1/aes_core/SB1/n2625 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U320  ( .A0(\U1/aes_core/SB1/n2826 ), 
        .A1(\U1/aes_core/SB1/n2866 ), .B0(\U1/aes_core/SB1/n2941 ), .Y(
        \U1/aes_core/SB1/n2624 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U319  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2939 ), .Y(\U1/aes_core/SB1/n2793 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U318  ( .A(\U1/aes_core/SB1/n2626 ), .B(
        \U1/aes_core/SB1/n2625 ), .C(\U1/aes_core/SB1/n2624 ), .D(
        \U1/aes_core/SB1/n2793 ), .Y(\U1/aes_core/SB1/n2627 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U317  ( .A(\U1/aes_core/SB1/n2632 ), .B(
        \U1/aes_core/SB1/n2631 ), .C(\U1/aes_core/SB1/n2630 ), .D(
        \U1/aes_core/SB1/n2629 ), .E(\U1/aes_core/SB1/n2628 ), .F(
        \U1/aes_core/SB1/n2627 ), .Y(\U1/aes_core/SB1/n2962 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U316  ( .A0(\U1/aes_core/SB1/n2747 ), 
        .A1(\U1/aes_core/SB1/n2943 ), .B0(\U1/aes_core/SB1/n2951 ), .B1(
        \U1/aes_core/SB1/n2865 ), .C0(\U1/aes_core/SB1/n2962 ), .Y(
        \U1/aes_core/SB1/n2633 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U315  ( .A(\U1/aes_core/SB1/n2633 ), .Y(
        \U1/aes_core/SB1/n2640 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U314  ( .A(\U1/aes_core/SB1/n2874 ), .B(
        \U1/aes_core/SB1/n2661 ), .Y(\U1/aes_core/SB1/n2783 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U313  ( .A1N(\U1/aes_core/SB1/n2783 ), 
        .A0(\U1/aes_core/SB1/n2913 ), .B0(\U1/aes_core/SB1/n2864 ), .Y(
        \U1/aes_core/SB1/n2636 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U312  ( .A0(\U1/aes_core/SB1/n2832 ), 
        .A1(\U1/aes_core/SB1/n2740 ), .B0(\U1/aes_core/SB1/n2912 ), .Y(
        \U1/aes_core/SB1/n2635 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U311  ( .A0(\U1/aes_core/SB1/n2939 ), 
        .A1(\U1/aes_core/SB1/n2873 ), .B0(\U1/aes_core/SB1/n2933 ), .Y(
        \U1/aes_core/SB1/n2634 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U310  ( .A(\U1/aes_core/SB1/n2910 ), .B(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2690 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U309  ( .A(\U1/aes_core/SB1/n2636 ), .B(
        \U1/aes_core/SB1/n2635 ), .C(\U1/aes_core/SB1/n2634 ), .D(
        \U1/aes_core/SB1/n2690 ), .Y(\U1/aes_core/SB1/n2639 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U308  ( .A(\U1/aes_core/SB1/n2909 ), .B(
        \U1/aes_core/SB1/n2941 ), .Y(\U1/aes_core/SB1/n2940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U307  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2866 ), .Y(\U1/aes_core/SB1/n2637 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U306  ( .A0(\U1/aes_core/SB1/n2940 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2637 ), .B1(
        \U1/aes_core/SB1/n2921 ), .C0(\U1/aes_core/SB1/n2843 ), .C1(
        \U1/aes_core/SB1/n2845 ), .Y(\U1/aes_core/SB1/n2638 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U305  ( .A(\U1/aes_core/SB1/n2643 ), .B(
        \U1/aes_core/SB1/n2642 ), .C(\U1/aes_core/SB1/n2641 ), .D(
        \U1/aes_core/SB1/n2640 ), .E(\U1/aes_core/SB1/n2639 ), .F(
        \U1/aes_core/SB1/n2638 ), .Y(\U1/aes_core/sb1 [26]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U304  ( .A(\U1/aes_core/SB1/n2747 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2945 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U303  ( .AN(\U1/aes_core/SB1/n2646 ), 
        .B(\U1/aes_core/SB1/n2645 ), .C(\U1/aes_core/SB1/n2644 ), .D(
        \U1/aes_core/SB1/n2945 ), .Y(\U1/aes_core/SB1/n2653 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U302  ( .A0(\U1/aes_core/SB1/n2647 ), 
        .A1(\U1/aes_core/SB1/n2912 ), .B0(\U1/aes_core/SB1/n2809 ), .Y(
        \U1/aes_core/SB1/n2649 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U299  ( .A(\U1/aes_core/SB1/n2865 ), .B(
        \U1/aes_core/SB1/n2933 ), .Y(\U1/aes_core/SB1/n2876 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U298  ( .A0(\U1/aes_core/SB1/n2755 ), 
        .A1(\U1/aes_core/SB1/n2955 ), .B0(\U1/aes_core/SB1/n2876 ), .B1(
        \U1/aes_core/SB1/n2908 ), .C0(\U1/aes_core/SB1/n2949 ), .C1(
        \U1/aes_core/SB1/n2958 ), .Y(\U1/aes_core/SB1/n2651 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U297  ( .A(\U1/aes_core/SB1/n2656 ), .B(
        \U1/aes_core/SB1/n2655 ), .C(\U1/aes_core/SB1/n2654 ), .D(
        \U1/aes_core/SB1/n2653 ), .E(\U1/aes_core/SB1/n2652 ), .F(
        \U1/aes_core/SB1/n2651 ), .Y(\U1/aes_core/SB1/n2839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U296  ( .AN(\U1/aes_core/SB1/n2660 ), 
        .B(\U1/aes_core/SB1/n2659 ), .C(\U1/aes_core/SB1/n2658 ), .D(
        \U1/aes_core/SB1/n2657 ), .Y(\U1/aes_core/SB1/n2670 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U295  ( .A0(\U1/aes_core/SB1/n2943 ), 
        .A1(\U1/aes_core/SB1/n2832 ), .B0(\U1/aes_core/SB1/n2938 ), .B1(
        \U1/aes_core/SB1/n2831 ), .C0(\U1/aes_core/SB1/n2661 ), .C1(
        \U1/aes_core/SB1/n2953 ), .Y(\U1/aes_core/SB1/n2669 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U294  ( .A0(\U1/aes_core/SB1/n2907 ), 
        .A1(\U1/aes_core/SB1/n2792 ), .B0(\U1/aes_core/SB1/n2662 ), .B1(
        \U1/aes_core/SB1/n2755 ), .Y(\U1/aes_core/SB1/n2663 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U293  ( .A0(\U1/aes_core/SB1/n2809 ), 
        .A1(\U1/aes_core/SB1/n2826 ), .B0(\U1/aes_core/SB1/n2825 ), .B1(
        \U1/aes_core/SB1/n2910 ), .C0(\U1/aes_core/SB1/n2663 ), .Y(
        \U1/aes_core/SB1/n2668 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U292  ( .A(\U1/aes_core/SB1/n2918 ), .B(
        \U1/aes_core/SB1/n2957 ), .Y(\U1/aes_core/SB1/n2665 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U291  ( .A0(\U1/aes_core/SB1/n2747 ), 
        .A1(\U1/aes_core/SB1/n2666 ), .B0(\U1/aes_core/SB1/n2939 ), .B1(
        \U1/aes_core/SB1/n2665 ), .C0(\U1/aes_core/SB1/n2664 ), .Y(
        \U1/aes_core/SB1/n2667 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U290  ( .AN(\U1/aes_core/SB1/n2670 ), 
        .B(\U1/aes_core/SB1/n2669 ), .C(\U1/aes_core/SB1/n2668 ), .D(
        \U1/aes_core/SB1/n2667 ), .Y(\U1/aes_core/SB1/n2884 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U289  ( .A(\U1/aes_core/SB1/n2671 ), .Y(
        \U1/aes_core/SB1/n2687 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U288  ( .A0(\U1/aes_core/SB1/n2776 ), 
        .A1(\U1/aes_core/SB1/n2845 ), .B0(\U1/aes_core/SB1/n2672 ), .Y(
        \U1/aes_core/SB1/n2686 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U287  ( .A0(\U1/aes_core/SB1/n2939 ), 
        .A1(\U1/aes_core/SB1/n2938 ), .B0(\U1/aes_core/SB1/n2909 ), .B1(
        \U1/aes_core/SB1/n2673 ), .Y(\U1/aes_core/SB1/n2674 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U286  ( .A0(\U1/aes_core/SB1/n2920 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2936 ), .B1(
        \U1/aes_core/SB1/n2948 ), .C0(\U1/aes_core/SB1/n2674 ), .Y(
        \U1/aes_core/SB1/n2685 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U285  ( .A(\U1/aes_core/SB1/n2678 ), .B(
        \U1/aes_core/SB1/n2677 ), .C(\U1/aes_core/SB1/n2676 ), .D(
        \U1/aes_core/SB1/n2675 ), .Y(\U1/aes_core/SB1/n2684 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U284  ( .AN(\U1/aes_core/SB1/n2682 ), 
        .B(\U1/aes_core/SB1/n2681 ), .C(\U1/aes_core/SB1/n2680 ), .D(
        \U1/aes_core/SB1/n2679 ), .Y(\U1/aes_core/SB1/n2683 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U283  ( .A(\U1/aes_core/SB1/n2688 ), .B(
        \U1/aes_core/SB1/n2687 ), .C(\U1/aes_core/SB1/n2686 ), .D(
        \U1/aes_core/SB1/n2685 ), .E(\U1/aes_core/SB1/n2684 ), .F(
        \U1/aes_core/SB1/n2683 ), .Y(\U1/aes_core/SB1/n2788 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U282  ( .A0(\U1/aes_core/SB1/n2875 ), 
        .A1(\U1/aes_core/SB1/n2792 ), .B0(\U1/aes_core/SB1/n2689 ), .Y(
        \U1/aes_core/SB1/n2704 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U281  ( .AN(\U1/aes_core/SB1/n2693 ), 
        .B(\U1/aes_core/SB1/n2692 ), .C(\U1/aes_core/SB1/n2691 ), .D(
        \U1/aes_core/SB1/n2690 ), .Y(\U1/aes_core/SB1/n2703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U280  ( .A(\U1/aes_core/SB1/n2930 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2944 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U279  ( .A(\U1/aes_core/SB1/n2696 ), .B(
        \U1/aes_core/SB1/n2695 ), .C(\U1/aes_core/SB1/n2694 ), .D(
        \U1/aes_core/SB1/n2944 ), .Y(\U1/aes_core/SB1/n2702 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U278  ( .A(\U1/aes_core/SB1/n2700 ), .B(
        \U1/aes_core/SB1/n2699 ), .C(\U1/aes_core/SB1/n2698 ), .D(
        \U1/aes_core/SB1/n2697 ), .Y(\U1/aes_core/SB1/n2701 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U277  ( .A(\U1/aes_core/SB1/n2706 ), .B(
        \U1/aes_core/SB1/n2705 ), .C(\U1/aes_core/SB1/n2704 ), .D(
        \U1/aes_core/SB1/n2703 ), .E(\U1/aes_core/SB1/n2702 ), .F(
        \U1/aes_core/SB1/n2701 ), .Y(\U1/aes_core/SB1/n2812 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U276  ( .AN(\U1/aes_core/SB1/n2710 ), 
        .B(\U1/aes_core/SB1/n2709 ), .C(\U1/aes_core/SB1/n2708 ), .D(
        \U1/aes_core/SB1/n2707 ), .Y(\U1/aes_core/SB1/n2719 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U275  ( .A(\U1/aes_core/SB1/n2714 ), .B(
        \U1/aes_core/SB1/n2713 ), .C(\U1/aes_core/SB1/n2712 ), .D(
        \U1/aes_core/SB1/n2711 ), .Y(\U1/aes_core/SB1/n2718 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U274  ( .A(\U1/aes_core/SB1/n2874 ), .B(
        \U1/aes_core/SB1/n2931 ), .C(\U1/aes_core/SB1/n2933 ), .Y(
        \U1/aes_core/SB1/n2716 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U273  ( .A0(\U1/aes_core/SB1/n2716 ), 
        .A1(\U1/aes_core/SB1/n2921 ), .B0(\U1/aes_core/SB1/n2755 ), .B1(
        \U1/aes_core/SB1/n2957 ), .C0(\U1/aes_core/SB1/n2715 ), .Y(
        \U1/aes_core/SB1/n2717 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U272  ( .A(\U1/aes_core/SB1/n2722 ), .B(
        \U1/aes_core/SB1/n2721 ), .C(\U1/aes_core/SB1/n2720 ), .D(
        \U1/aes_core/SB1/n2719 ), .E(\U1/aes_core/SB1/n2718 ), .F(
        \U1/aes_core/SB1/n2717 ), .Y(\U1/aes_core/SB1/n2860 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U271  ( .A0(\U1/aes_core/SB1/n2755 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2723 ), .Y(
        \U1/aes_core/SB1/n2737 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U270  ( .A0(\U1/aes_core/SB1/n2864 ), 
        .A1(\U1/aes_core/SB1/n2866 ), .B0(\U1/aes_core/SB1/n2942 ), .B1(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2724 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U269  ( .A0(\U1/aes_core/SB1/n2775 ), 
        .A1(\U1/aes_core/SB1/n2863 ), .B0(\U1/aes_core/SB1/n2776 ), .B1(
        \U1/aes_core/SB1/n2840 ), .C0(\U1/aes_core/SB1/n2724 ), .Y(
        \U1/aes_core/SB1/n2736 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U268  ( .A(\U1/aes_core/SB1/n2725 ), .Y(
        \U1/aes_core/SB1/n2728 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U267  ( .AN(\U1/aes_core/SB1/n2729 ), 
        .B(\U1/aes_core/SB1/n2728 ), .C(\U1/aes_core/SB1/n2727 ), .D(
        \U1/aes_core/SB1/n2726 ), .Y(\U1/aes_core/SB1/n2735 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U266  ( .A(\U1/aes_core/SB1/n2733 ), .B(
        \U1/aes_core/SB1/n2732 ), .C(\U1/aes_core/SB1/n2731 ), .D(
        \U1/aes_core/SB1/n2730 ), .Y(\U1/aes_core/SB1/n2734 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U265  ( .A(\U1/aes_core/SB1/n2739 ), .B(
        \U1/aes_core/SB1/n2738 ), .C(\U1/aes_core/SB1/n2737 ), .D(
        \U1/aes_core/SB1/n2736 ), .E(\U1/aes_core/SB1/n2735 ), .F(
        \U1/aes_core/SB1/n2734 ), .Y(\U1/aes_core/SB1/n2819 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U264  ( .A0(\U1/aes_core/SB1/n2931 ), 
        .A1(\U1/aes_core/SB1/n2740 ), .B0(\U1/aes_core/SB1/n2941 ), .B1(
        \U1/aes_core/SB1/n2866 ), .Y(\U1/aes_core/SB1/n2741 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U263  ( .A0(\U1/aes_core/SB1/n2792 ), 
        .A1(\U1/aes_core/SB1/n2958 ), .B0(\U1/aes_core/SB1/n2742 ), .B1(
        \U1/aes_core/SB1/n2948 ), .C0(\U1/aes_core/SB1/n2741 ), .Y(
        \U1/aes_core/SB1/n2754 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U262  ( .AN(\U1/aes_core/SB1/n2746 ), 
        .B(\U1/aes_core/SB1/n2745 ), .C(\U1/aes_core/SB1/n2744 ), .D(
        \U1/aes_core/SB1/n2743 ), .Y(\U1/aes_core/SB1/n2753 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U261  ( .A0(\U1/aes_core/SB1/n2951 ), 
        .A1(\U1/aes_core/SB1/n2747 ), .B0(\U1/aes_core/SB1/n2942 ), .Y(
        \U1/aes_core/SB1/n2751 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U260  ( .A(\U1/aes_core/SB1/n2918 ), .B(
        \U1/aes_core/SB1/n2923 ), .Y(\U1/aes_core/SB1/n2748 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U259  ( .A0(\U1/aes_core/SB1/n2873 ), 
        .A1(\U1/aes_core/SB1/n2748 ), .B0(\U1/aes_core/SB1/n2874 ), .B1(
        \U1/aes_core/SB1/n2820 ), .Y(\U1/aes_core/SB1/n2749 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U258  ( .A(\U1/aes_core/SB1/n2751 ), .B(
        \U1/aes_core/SB1/n2750 ), .C(\U1/aes_core/SB1/n2749 ), .Y(
        \U1/aes_core/SB1/n2752 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U257  ( .A(\U1/aes_core/SB1/n2812 ), .B(
        \U1/aes_core/SB1/n2860 ), .C(\U1/aes_core/SB1/n2819 ), .D(
        \U1/aes_core/SB1/n2754 ), .E(\U1/aes_core/SB1/n2753 ), .F(
        \U1/aes_core/SB1/n2752 ), .Y(\U1/aes_core/SB1/n2927 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U256  ( .A(\U1/aes_core/SB1/n2839 ), .B(
        \U1/aes_core/SB1/n2884 ), .C(\U1/aes_core/SB1/n2788 ), .D(
        \U1/aes_core/SB1/n2927 ), .Y(\U1/aes_core/SB1/n2768 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U255  ( .A0(\U1/aes_core/SB1/n2907 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2755 ), .B1(
        \U1/aes_core/SB1/n2923 ), .Y(\U1/aes_core/SB1/n2756 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U254  ( .A0(\U1/aes_core/SB1/n2912 ), 
        .A1(\U1/aes_core/SB1/n2930 ), .B0(\U1/aes_core/SB1/n2943 ), .B1(
        \U1/aes_core/SB1/n2951 ), .C0(\U1/aes_core/SB1/n2756 ), .Y(
        \U1/aes_core/SB1/n2767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U253  ( .A(\U1/aes_core/SB1/n2757 ), .Y(
        \U1/aes_core/SB1/n2760 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U252  ( .A0(\U1/aes_core/SB1/n2758 ), 
        .A1(\U1/aes_core/SB1/n2863 ), .B0(\U1/aes_core/SB1/n2791 ), .B1(
        \U1/aes_core/SB1/n2843 ), .Y(\U1/aes_core/SB1/n2759 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U251  ( .A0(\U1/aes_core/SB1/n2931 ), 
        .A1(\U1/aes_core/SB1/n2760 ), .B0(\U1/aes_core/SB1/n2913 ), .B1(
        \U1/aes_core/SB1/n2841 ), .C0(\U1/aes_core/SB1/n2759 ), .Y(
        \U1/aes_core/SB1/n2766 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U250  ( .A0(\U1/aes_core/SB1/n2953 ), 
        .A1(\U1/aes_core/SB1/n2809 ), .B0(\U1/aes_core/SB1/n2933 ), .Y(
        \U1/aes_core/SB1/n2764 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB1/U249  ( .A(\U1/aes_core/SB1/n2764 ), .B(
        \U1/aes_core/SB1/n2763 ), .C(\U1/aes_core/SB1/n2762 ), .D(
        \U1/aes_core/SB1/n2761 ), .Y(\U1/aes_core/SB1/n2765 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U248  ( .AN(\U1/aes_core/SB1/n2768 ), 
        .B(\U1/aes_core/SB1/n2767 ), .C(\U1/aes_core/SB1/n2766 ), .D(
        \U1/aes_core/SB1/n2765 ), .Y(\U1/aes_core/sb1 [27]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U247  ( .A0(\U1/aes_core/SB1/n2783 ), 
        .A1(\U1/aes_core/SB1/n2919 ), .B0(\U1/aes_core/SB1/n2842 ), .Y(
        \U1/aes_core/SB1/n2780 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U246  ( .A(\U1/aes_core/SB1/n2771 ), .B(
        \U1/aes_core/SB1/n2770 ), .C(\U1/aes_core/SB1/n2769 ), .Y(
        \U1/aes_core/SB1/n2779 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U245  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2942 ), .Y(\U1/aes_core/SB1/n2774 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U244  ( .A(\U1/aes_core/SB1/n2913 ), .B(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2772 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U243  ( .A0(\U1/aes_core/SB1/n2774 ), 
        .A1(\U1/aes_core/SB1/n2773 ), .B0(\U1/aes_core/SB1/n2772 ), .B1(
        \U1/aes_core/SB1/n2936 ), .C0(\U1/aes_core/SB1/n2919 ), .C1(
        \U1/aes_core/SB1/n2824 ), .Y(\U1/aes_core/SB1/n2778 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U242  ( .A0(\U1/aes_core/SB1/n2875 ), 
        .A1(\U1/aes_core/SB1/n2776 ), .B0(\U1/aes_core/SB1/n2958 ), .B1(
        \U1/aes_core/SB1/n2948 ), .C0(\U1/aes_core/SB1/n2921 ), .C1(
        \U1/aes_core/SB1/n2775 ), .Y(\U1/aes_core/SB1/n2777 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U241  ( .A(\U1/aes_core/SB1/n2782 ), .B(
        \U1/aes_core/SB1/n2781 ), .C(\U1/aes_core/SB1/n2780 ), .D(
        \U1/aes_core/SB1/n2779 ), .E(\U1/aes_core/SB1/n2778 ), .F(
        \U1/aes_core/SB1/n2777 ), .Y(\U1/aes_core/SB1/n2928 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U240  ( .A0(\U1/aes_core/SB1/n2783 ), 
        .A1(\U1/aes_core/SB1/n2792 ), .B0(\U1/aes_core/SB1/n2863 ), .Y(
        \U1/aes_core/SB1/n2818 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB1/U239  ( .A0(\U1/aes_core/SB1/n2908 ), 
        .A1(\U1/aes_core/SB1/n2921 ), .A2(\U1/aes_core/SB1/n2840 ), .B0(
        \U1/aes_core/SB1/n2937 ), .Y(\U1/aes_core/SB1/n2817 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U238  ( .A(\U1/aes_core/SB1/n2787 ), .B(
        \U1/aes_core/SB1/n2786 ), .C(\U1/aes_core/SB1/n2785 ), .D(
        \U1/aes_core/SB1/n2784 ), .Y(\U1/aes_core/SB1/n2814 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U237  ( .A(\U1/aes_core/SB1/n2788 ), .Y(
        \U1/aes_core/SB1/n2811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U236  ( .A(\U1/aes_core/SB1/n2789 ), .Y(
        \U1/aes_core/SB1/n2805 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB1/U235  ( .A0(\U1/aes_core/SB1/n2791 ), 
        .A1(\U1/aes_core/SB1/n2949 ), .B0N(\U1/aes_core/SB1/n2790 ), .Y(
        \U1/aes_core/SB1/n2804 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U234  ( .A0(\U1/aes_core/SB1/n2956 ), 
        .A1(\U1/aes_core/SB1/n2792 ), .B0(\U1/aes_core/SB1/n2842 ), .B1(
        \U1/aes_core/SB1/n2923 ), .C0(\U1/aes_core/SB1/n2937 ), .C1(
        \U1/aes_core/SB1/n2958 ), .Y(\U1/aes_core/SB1/n2803 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U233  ( .AN(\U1/aes_core/SB1/n2796 ), 
        .B(\U1/aes_core/SB1/n2795 ), .C(\U1/aes_core/SB1/n2794 ), .D(
        \U1/aes_core/SB1/n2793 ), .Y(\U1/aes_core/SB1/n2802 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U232  ( .A(\U1/aes_core/SB1/n2800 ), .B(
        \U1/aes_core/SB1/n2799 ), .C(\U1/aes_core/SB1/n2798 ), .D(
        \U1/aes_core/SB1/n2797 ), .Y(\U1/aes_core/SB1/n2801 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U231  ( .A(\U1/aes_core/SB1/n2806 ), .B(
        \U1/aes_core/SB1/n2805 ), .C(\U1/aes_core/SB1/n2804 ), .D(
        \U1/aes_core/SB1/n2803 ), .E(\U1/aes_core/SB1/n2802 ), .F(
        \U1/aes_core/SB1/n2801 ), .Y(\U1/aes_core/SB1/n2807 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U230  ( .A(\U1/aes_core/SB1/n2807 ), .Y(
        \U1/aes_core/SB1/n2906 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U229  ( .A0(\U1/aes_core/SB1/n2875 ), 
        .A1(\U1/aes_core/SB1/n2918 ), .B0(\U1/aes_core/SB1/n2958 ), .B1(
        \U1/aes_core/SB1/n2957 ), .Y(\U1/aes_core/SB1/n2808 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U228  ( .A0(\U1/aes_core/SB1/n2865 ), 
        .A1(\U1/aes_core/SB1/n2809 ), .B0(\U1/aes_core/SB1/n2910 ), .B1(
        \U1/aes_core/SB1/n2932 ), .C0(\U1/aes_core/SB1/n2808 ), .Y(
        \U1/aes_core/SB1/n2810 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U227  ( .AN(\U1/aes_core/SB1/n2812 ), 
        .B(\U1/aes_core/SB1/n2811 ), .C(\U1/aes_core/SB1/n2906 ), .D(
        \U1/aes_core/SB1/n2810 ), .Y(\U1/aes_core/SB1/n2813 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U226  ( .A(\U1/aes_core/SB1/n2818 ), .B(
        \U1/aes_core/SB1/n2817 ), .C(\U1/aes_core/SB1/n2816 ), .D(
        \U1/aes_core/SB1/n2815 ), .E(\U1/aes_core/SB1/n2814 ), .F(
        \U1/aes_core/SB1/n2813 ), .Y(\U1/aes_core/SB1/n2883 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U225  ( .A(\U1/aes_core/SB1/n2819 ), .Y(
        \U1/aes_core/SB1/n2823 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U224  ( .A0(\U1/aes_core/SB1/n2821 ), 
        .A1(\U1/aes_core/SB1/n2820 ), .B0(\U1/aes_core/SB1/n2867 ), .B1(
        \U1/aes_core/SB1/n2826 ), .Y(\U1/aes_core/SB1/n2822 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U223  ( .A0(\U1/aes_core/SB1/n2937 ), 
        .A1(\U1/aes_core/SB1/n2824 ), .B0(\U1/aes_core/SB1/n2823 ), .C0(
        \U1/aes_core/SB1/n2822 ), .Y(\U1/aes_core/SB1/n2838 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U222  ( .A0(\U1/aes_core/SB1/n2825 ), 
        .A1(\U1/aes_core/SB1/n2909 ), .B0(\U1/aes_core/SB1/n2938 ), .Y(
        \U1/aes_core/SB1/n2830 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U221  ( .A0(\U1/aes_core/SB1/n2826 ), 
        .A1(\U1/aes_core/SB1/n2912 ), .B0(\U1/aes_core/SB1/n2941 ), .Y(
        \U1/aes_core/SB1/n2829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U220  ( .A(\U1/aes_core/SB1/n2830 ), .B(
        \U1/aes_core/SB1/n2829 ), .C(\U1/aes_core/SB1/n2828 ), .D(
        \U1/aes_core/SB1/n2827 ), .Y(\U1/aes_core/SB1/n2837 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U219  ( .A(\U1/aes_core/SB1/n2868 ), .B(
        \U1/aes_core/SB1/n2831 ), .Y(\U1/aes_core/SB1/n2835 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U218  ( .A(\U1/aes_core/SB1/n2832 ), .B(
        \U1/aes_core/SB1/n2873 ), .Y(\U1/aes_core/SB1/n2834 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U217  ( .A0(\U1/aes_core/SB1/n2835 ), 
        .A1(\U1/aes_core/SB1/n2955 ), .B0(\U1/aes_core/SB1/n2834 ), .B1(
        \U1/aes_core/SB1/n2919 ), .C0(\U1/aes_core/SB1/n2833 ), .C1(
        \U1/aes_core/SB1/n2920 ), .Y(\U1/aes_core/SB1/n2836 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U216  ( .A(\U1/aes_core/SB1/n2928 ), .B(
        \U1/aes_core/SB1/n2883 ), .C(\U1/aes_core/SB1/n2839 ), .D(
        \U1/aes_core/SB1/n2838 ), .E(\U1/aes_core/SB1/n2837 ), .F(
        \U1/aes_core/SB1/n2836 ), .Y(\U1/aes_core/sb1 [28]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U215  ( .A1N(\U1/aes_core/SB1/n2841 ), 
        .A0(\U1/aes_core/SB1/n2840 ), .B0(\U1/aes_core/SB1/n2918 ), .Y(
        \U1/aes_core/SB1/n2857 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U214  ( .A(\U1/aes_core/SB1/n2931 ), .B(
        \U1/aes_core/SB1/n2912 ), .Y(\U1/aes_core/SB1/n2844 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U213  ( .A0(\U1/aes_core/SB1/n2955 ), 
        .A1(\U1/aes_core/SB1/n2845 ), .B0(\U1/aes_core/SB1/n2844 ), .B1(
        \U1/aes_core/SB1/n2958 ), .C0(\U1/aes_core/SB1/n2843 ), .C1(
        \U1/aes_core/SB1/n2842 ), .Y(\U1/aes_core/SB1/n2856 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U212  ( .A(\U1/aes_core/SB1/n2846 ), .Y(
        \U1/aes_core/SB1/n2849 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U211  ( .AN(\U1/aes_core/SB1/n2850 ), 
        .B(\U1/aes_core/SB1/n2849 ), .C(\U1/aes_core/SB1/n2848 ), .D(
        \U1/aes_core/SB1/n2847 ), .Y(\U1/aes_core/SB1/n2855 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U210  ( .A(\U1/aes_core/SB1/n2853 ), .B(
        \U1/aes_core/SB1/n2852 ), .C(\U1/aes_core/SB1/n2851 ), .Y(
        \U1/aes_core/SB1/n2854 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U209  ( .A(\U1/aes_core/SB1/n2859 ), .B(
        \U1/aes_core/SB1/n2858 ), .C(\U1/aes_core/SB1/n2857 ), .D(
        \U1/aes_core/SB1/n2856 ), .E(\U1/aes_core/SB1/n2855 ), .F(
        \U1/aes_core/SB1/n2854 ), .Y(\U1/aes_core/SB1/n2929 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U208  ( .A(\U1/aes_core/SB1/n2860 ), .Y(
        \U1/aes_core/SB1/n2862 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U207  ( .A0(\U1/aes_core/SB1/n2942 ), 
        .A1(\U1/aes_core/SB1/n2939 ), .B0(\U1/aes_core/SB1/n2943 ), .B1(
        \U1/aes_core/SB1/n2941 ), .Y(\U1/aes_core/SB1/n2861 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U206  ( .A0(\U1/aes_core/SB1/n2918 ), 
        .A1(\U1/aes_core/SB1/n2863 ), .B0(\U1/aes_core/SB1/n2862 ), .C0(
        \U1/aes_core/SB1/n2861 ), .Y(\U1/aes_core/SB1/n2882 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U205  ( .A0(\U1/aes_core/SB1/n2865 ), 
        .A1(\U1/aes_core/SB1/n2942 ), .B0(\U1/aes_core/SB1/n2864 ), .Y(
        \U1/aes_core/SB1/n2871 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U204  ( .A0(\U1/aes_core/SB1/n2868 ), 
        .A1(\U1/aes_core/SB1/n2867 ), .B0(\U1/aes_core/SB1/n2866 ), .Y(
        \U1/aes_core/SB1/n2870 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U203  ( .AN(\U1/aes_core/SB1/n2872 ), 
        .B(\U1/aes_core/SB1/n2871 ), .C(\U1/aes_core/SB1/n2870 ), .D(
        \U1/aes_core/SB1/n2869 ), .Y(\U1/aes_core/SB1/n2881 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U202  ( .A0(\U1/aes_core/SB1/n2938 ), 
        .A1(\U1/aes_core/SB1/n2874 ), .B0(\U1/aes_core/SB1/n2873 ), .Y(
        \U1/aes_core/SB1/n2878 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB1/U201  ( .A0(\U1/aes_core/SB1/n2920 ), .A1(
        \U1/aes_core/SB1/n2876 ), .B0(\U1/aes_core/SB1/n2957 ), .B1(
        \U1/aes_core/SB1/n2875 ), .Y(\U1/aes_core/SB1/n2877 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U200  ( .A0(\U1/aes_core/SB1/n2879 ), 
        .A1(\U1/aes_core/SB1/n2919 ), .B0(\U1/aes_core/SB1/n2878 ), .C0(
        \U1/aes_core/SB1/n2877 ), .Y(\U1/aes_core/SB1/n2880 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U199  ( .A(\U1/aes_core/SB1/n2929 ), .B(
        \U1/aes_core/SB1/n2884 ), .C(\U1/aes_core/SB1/n2883 ), .D(
        \U1/aes_core/SB1/n2882 ), .E(\U1/aes_core/SB1/n2881 ), .F(
        \U1/aes_core/SB1/n2880 ), .Y(\U1/aes_core/sb1 [29]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U198  ( .A0(\U1/aes_core/SB1/n3212 ), 
        .A1(\U1/aes_core/SB1/n3232 ), .B0(\U1/aes_core/SB1/n3253 ), .B1(
        \U1/aes_core/SB1/n3243 ), .Y(\U1/aes_core/SB1/n2885 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U197  ( .A0(\U1/aes_core/SB1/n3163 ), 
        .A1(\U1/aes_core/SB1/n3257 ), .B0(\U1/aes_core/SB1/n3113 ), .B1(
        \U1/aes_core/SB1/n3184 ), .C0(\U1/aes_core/SB1/n2885 ), .Y(
        \U1/aes_core/SB1/n2891 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U196  ( .A(\U1/aes_core/SB1/n3238 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3047 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U195  ( .A(\U1/aes_core/SB1/n3212 ), .B(
        \U1/aes_core/SB1/n3188 ), .Y(\U1/aes_core/SB1/n3028 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U194  ( .A(\U1/aes_core/SB1/n3232 ), .B(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n2996 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U193  ( .A(\U1/aes_core/SB1/n3152 ), .B(
        \U1/aes_core/SB1/n3195 ), .Y(\U1/aes_core/SB1/n3015 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U192  ( .A(\U1/aes_core/SB1/n3047 ), .B(
        \U1/aes_core/SB1/n3028 ), .C(\U1/aes_core/SB1/n2996 ), .D(
        \U1/aes_core/SB1/n3015 ), .Y(\U1/aes_core/SB1/n2890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U191  ( .A(\U1/aes_core/SB1/n3258 ), .B(
        \U1/aes_core/SB1/n3236 ), .Y(\U1/aes_core/SB1/n3141 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U190  ( .A0(\U1/aes_core/SB1/n3189 ), 
        .A1(\U1/aes_core/SB1/n3141 ), .B0(\U1/aes_core/SB1/n3242 ), .Y(
        \U1/aes_core/SB1/n2888 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U189  ( .A0(\U1/aes_core/SB1/n3239 ), 
        .A1(\U1/aes_core/SB1/n3130 ), .B0(\U1/aes_core/SB1/n3142 ), .Y(
        \U1/aes_core/SB1/n2887 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U188  ( .A0(\U1/aes_core/SB1/n3147 ), 
        .A1(\U1/aes_core/SB1/n3187 ), .B0(\U1/aes_core/SB1/n3241 ), .Y(
        \U1/aes_core/SB1/n2886 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U187  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3239 ), .Y(\U1/aes_core/SB1/n3114 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U186  ( .A(\U1/aes_core/SB1/n2888 ), .B(
        \U1/aes_core/SB1/n2887 ), .C(\U1/aes_core/SB1/n2886 ), .D(
        \U1/aes_core/SB1/n3114 ), .Y(\U1/aes_core/SB1/n2889 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U185  ( .A(\U1/aes_core/SB1/n2894 ), .B(
        \U1/aes_core/SB1/n2893 ), .C(\U1/aes_core/SB1/n2892 ), .D(
        \U1/aes_core/SB1/n2891 ), .E(\U1/aes_core/SB1/n2890 ), .F(
        \U1/aes_core/SB1/n2889 ), .Y(\U1/aes_core/SB1/n3262 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U184  ( .A0(\U1/aes_core/SB1/n3068 ), 
        .A1(\U1/aes_core/SB1/n3243 ), .B0(\U1/aes_core/SB1/n3251 ), .B1(
        \U1/aes_core/SB1/n3186 ), .C0(\U1/aes_core/SB1/n3262 ), .Y(
        \U1/aes_core/SB1/n2895 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U183  ( .A(\U1/aes_core/SB1/n2895 ), .Y(
        \U1/aes_core/SB1/n2902 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U182  ( .A(\U1/aes_core/SB1/n3195 ), .B(
        \U1/aes_core/SB1/n2982 ), .Y(\U1/aes_core/SB1/n3104 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U181  ( .A1N(\U1/aes_core/SB1/n3104 ), 
        .A0(\U1/aes_core/SB1/n3213 ), .B0(\U1/aes_core/SB1/n3185 ), .Y(
        \U1/aes_core/SB1/n2898 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U180  ( .A0(\U1/aes_core/SB1/n3153 ), 
        .A1(\U1/aes_core/SB1/n3061 ), .B0(\U1/aes_core/SB1/n3212 ), .Y(
        \U1/aes_core/SB1/n2897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U179  ( .A0(\U1/aes_core/SB1/n3239 ), 
        .A1(\U1/aes_core/SB1/n3194 ), .B0(\U1/aes_core/SB1/n3233 ), .Y(
        \U1/aes_core/SB1/n2896 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U178  ( .A(\U1/aes_core/SB1/n3210 ), .B(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n3011 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U177  ( .A(\U1/aes_core/SB1/n2898 ), .B(
        \U1/aes_core/SB1/n2897 ), .C(\U1/aes_core/SB1/n2896 ), .D(
        \U1/aes_core/SB1/n3011 ), .Y(\U1/aes_core/SB1/n2901 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U176  ( .A(\U1/aes_core/SB1/n3209 ), .B(
        \U1/aes_core/SB1/n3241 ), .Y(\U1/aes_core/SB1/n3240 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U175  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3187 ), .Y(\U1/aes_core/SB1/n2899 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U174  ( .A0(\U1/aes_core/SB1/n3240 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n2899 ), .B1(
        \U1/aes_core/SB1/n3221 ), .C0(\U1/aes_core/SB1/n3164 ), .C1(
        \U1/aes_core/SB1/n3166 ), .Y(\U1/aes_core/SB1/n2900 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U173  ( .A(\U1/aes_core/SB1/n2905 ), .B(
        \U1/aes_core/SB1/n2904 ), .C(\U1/aes_core/SB1/n2903 ), .D(
        \U1/aes_core/SB1/n2902 ), .E(\U1/aes_core/SB1/n2901 ), .F(
        \U1/aes_core/SB1/n2900 ), .Y(\U1/aes_core/sb1 [2]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U172  ( .A0(\U1/aes_core/SB1/n2908 ), 
        .A1(\U1/aes_core/SB1/n2948 ), .B0(\U1/aes_core/SB1/n2907 ), .B1(
        \U1/aes_core/SB1/n2955 ), .C0(\U1/aes_core/SB1/n2906 ), .Y(
        \U1/aes_core/SB1/n2926 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U171  ( .A0(\U1/aes_core/SB1/n2909 ), 
        .A1(\U1/aes_core/SB1/n2953 ), .B0(\U1/aes_core/SB1/n2942 ), .Y(
        \U1/aes_core/SB1/n2917 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U170  ( .A0(\U1/aes_core/SB1/n2933 ), 
        .A1(\U1/aes_core/SB1/n2910 ), .B0(\U1/aes_core/SB1/n2941 ), .Y(
        \U1/aes_core/SB1/n2916 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U169  ( .A0(\U1/aes_core/SB1/n2913 ), 
        .A1(\U1/aes_core/SB1/n2912 ), .B0(\U1/aes_core/SB1/n2911 ), .Y(
        \U1/aes_core/SB1/n2915 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U168  ( .A(\U1/aes_core/SB1/n2917 ), .B(
        \U1/aes_core/SB1/n2916 ), .C(\U1/aes_core/SB1/n2915 ), .D(
        \U1/aes_core/SB1/n2914 ), .Y(\U1/aes_core/SB1/n2925 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U167  ( .A(\U1/aes_core/SB1/n2948 ), .B(
        \U1/aes_core/SB1/n2918 ), .Y(\U1/aes_core/SB1/n2950 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U166  ( .A(\U1/aes_core/SB1/n2938 ), .B(
        \U1/aes_core/SB1/n2950 ), .Y(\U1/aes_core/SB1/n2922 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U165  ( .A0(\U1/aes_core/SB1/n2936 ), 
        .A1(\U1/aes_core/SB1/n2923 ), .B0(\U1/aes_core/SB1/n2922 ), .B1(
        \U1/aes_core/SB1/n2921 ), .C0(\U1/aes_core/SB1/n2920 ), .C1(
        \U1/aes_core/SB1/n2919 ), .Y(\U1/aes_core/SB1/n2924 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U164  ( .A(\U1/aes_core/SB1/n2929 ), .B(
        \U1/aes_core/SB1/n2928 ), .C(\U1/aes_core/SB1/n2927 ), .D(
        \U1/aes_core/SB1/n2926 ), .E(\U1/aes_core/SB1/n2925 ), .F(
        \U1/aes_core/SB1/n2924 ), .Y(\U1/aes_core/sb1 [30]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U163  ( .A0(\U1/aes_core/SB1/n2933 ), 
        .A1(\U1/aes_core/SB1/n2932 ), .B0(\U1/aes_core/SB1/n2931 ), .B1(
        \U1/aes_core/SB1/n2930 ), .Y(\U1/aes_core/SB1/n2934 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U162  ( .A0(\U1/aes_core/SB1/n2937 ), 
        .A1(\U1/aes_core/SB1/n2936 ), .B0(\U1/aes_core/SB1/n2935 ), .C0(
        \U1/aes_core/SB1/n2934 ), .Y(\U1/aes_core/SB1/n2961 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U161  ( .A1N(\U1/aes_core/SB1/n2940 ), 
        .A0(\U1/aes_core/SB1/n2939 ), .B0(\U1/aes_core/SB1/n2938 ), .Y(
        \U1/aes_core/SB1/n2947 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U160  ( .A0(\U1/aes_core/SB1/n2943 ), 
        .A1(\U1/aes_core/SB1/n2942 ), .B0(\U1/aes_core/SB1/n2941 ), .Y(
        \U1/aes_core/SB1/n2946 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U159  ( .A(\U1/aes_core/SB1/n2947 ), .B(
        \U1/aes_core/SB1/n2946 ), .C(\U1/aes_core/SB1/n2945 ), .D(
        \U1/aes_core/SB1/n2944 ), .Y(\U1/aes_core/SB1/n2960 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U158  ( .A(\U1/aes_core/SB1/n2949 ), .B(
        \U1/aes_core/SB1/n2948 ), .Y(\U1/aes_core/SB1/n2952 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U157  ( .A0(\U1/aes_core/SB1/n2953 ), 
        .A1(\U1/aes_core/SB1/n2952 ), .B0(\U1/aes_core/SB1/n2951 ), .B1(
        \U1/aes_core/SB1/n2950 ), .Y(\U1/aes_core/SB1/n2954 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U156  ( .A0(\U1/aes_core/SB1/n2958 ), 
        .A1(\U1/aes_core/SB1/n2957 ), .B0(\U1/aes_core/SB1/n2956 ), .B1(
        \U1/aes_core/SB1/n2955 ), .C0(\U1/aes_core/SB1/n2954 ), .Y(
        \U1/aes_core/SB1/n2959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U155  ( .A(\U1/aes_core/SB1/n2964 ), .B(
        \U1/aes_core/SB1/n2963 ), .C(\U1/aes_core/SB1/n2962 ), .D(
        \U1/aes_core/SB1/n2961 ), .E(\U1/aes_core/SB1/n2960 ), .F(
        \U1/aes_core/SB1/n2959 ), .Y(\U1/aes_core/sb1 [31]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U154  ( .A(\U1/aes_core/SB1/n3068 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3245 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U153  ( .AN(\U1/aes_core/SB1/n2967 ), 
        .B(\U1/aes_core/SB1/n2966 ), .C(\U1/aes_core/SB1/n2965 ), .D(
        \U1/aes_core/SB1/n3245 ), .Y(\U1/aes_core/SB1/n2974 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U152  ( .A0(\U1/aes_core/SB1/n2968 ), 
        .A1(\U1/aes_core/SB1/n3212 ), .B0(\U1/aes_core/SB1/n3130 ), .Y(
        \U1/aes_core/SB1/n2970 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U149  ( .A(\U1/aes_core/SB1/n3186 ), .B(
        \U1/aes_core/SB1/n3233 ), .Y(\U1/aes_core/SB1/n3197 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U148  ( .A0(\U1/aes_core/SB1/n3076 ), 
        .A1(\U1/aes_core/SB1/n3255 ), .B0(\U1/aes_core/SB1/n3197 ), .B1(
        \U1/aes_core/SB1/n3208 ), .C0(\U1/aes_core/SB1/n3249 ), .C1(
        \U1/aes_core/SB1/n3258 ), .Y(\U1/aes_core/SB1/n2972 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U147  ( .A(\U1/aes_core/SB1/n2977 ), .B(
        \U1/aes_core/SB1/n2976 ), .C(\U1/aes_core/SB1/n2975 ), .D(
        \U1/aes_core/SB1/n2974 ), .E(\U1/aes_core/SB1/n2973 ), .F(
        \U1/aes_core/SB1/n2972 ), .Y(\U1/aes_core/SB1/n3160 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U146  ( .AN(\U1/aes_core/SB1/n2981 ), 
        .B(\U1/aes_core/SB1/n2980 ), .C(\U1/aes_core/SB1/n2979 ), .D(
        \U1/aes_core/SB1/n2978 ), .Y(\U1/aes_core/SB1/n2991 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB1/U145  ( .A0(\U1/aes_core/SB1/n3243 ), 
        .A1(\U1/aes_core/SB1/n3153 ), .B0(\U1/aes_core/SB1/n3238 ), .B1(
        \U1/aes_core/SB1/n3152 ), .C0(\U1/aes_core/SB1/n2982 ), .C1(
        \U1/aes_core/SB1/n3253 ), .Y(\U1/aes_core/SB1/n2990 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U144  ( .A0(\U1/aes_core/SB1/n3207 ), 
        .A1(\U1/aes_core/SB1/n3113 ), .B0(\U1/aes_core/SB1/n2983 ), .B1(
        \U1/aes_core/SB1/n3076 ), .Y(\U1/aes_core/SB1/n2984 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U143  ( .A0(\U1/aes_core/SB1/n3130 ), 
        .A1(\U1/aes_core/SB1/n3147 ), .B0(\U1/aes_core/SB1/n3146 ), .B1(
        \U1/aes_core/SB1/n3210 ), .C0(\U1/aes_core/SB1/n2984 ), .Y(
        \U1/aes_core/SB1/n2989 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U142  ( .A(\U1/aes_core/SB1/n3218 ), .B(
        \U1/aes_core/SB1/n3257 ), .Y(\U1/aes_core/SB1/n2986 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U141  ( .A0(\U1/aes_core/SB1/n3068 ), 
        .A1(\U1/aes_core/SB1/n2987 ), .B0(\U1/aes_core/SB1/n3239 ), .B1(
        \U1/aes_core/SB1/n2986 ), .C0(\U1/aes_core/SB1/n2985 ), .Y(
        \U1/aes_core/SB1/n2988 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U140  ( .AN(\U1/aes_core/SB1/n2991 ), 
        .B(\U1/aes_core/SB1/n2990 ), .C(\U1/aes_core/SB1/n2989 ), .D(
        \U1/aes_core/SB1/n2988 ), .Y(\U1/aes_core/SB1/n3205 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U139  ( .A(\U1/aes_core/SB1/n2992 ), .Y(
        \U1/aes_core/SB1/n3008 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U138  ( .A0(\U1/aes_core/SB1/n3097 ), 
        .A1(\U1/aes_core/SB1/n3166 ), .B0(\U1/aes_core/SB1/n2993 ), .Y(
        \U1/aes_core/SB1/n3007 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U137  ( .A0(\U1/aes_core/SB1/n3239 ), 
        .A1(\U1/aes_core/SB1/n3238 ), .B0(\U1/aes_core/SB1/n3209 ), .B1(
        \U1/aes_core/SB1/n2994 ), .Y(\U1/aes_core/SB1/n2995 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U136  ( .A0(\U1/aes_core/SB1/n3220 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3236 ), .B1(
        \U1/aes_core/SB1/n3248 ), .C0(\U1/aes_core/SB1/n2995 ), .Y(
        \U1/aes_core/SB1/n3006 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U135  ( .A(\U1/aes_core/SB1/n2999 ), .B(
        \U1/aes_core/SB1/n2998 ), .C(\U1/aes_core/SB1/n2997 ), .D(
        \U1/aes_core/SB1/n2996 ), .Y(\U1/aes_core/SB1/n3005 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U134  ( .AN(\U1/aes_core/SB1/n3003 ), 
        .B(\U1/aes_core/SB1/n3002 ), .C(\U1/aes_core/SB1/n3001 ), .D(
        \U1/aes_core/SB1/n3000 ), .Y(\U1/aes_core/SB1/n3004 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U133  ( .A(\U1/aes_core/SB1/n3009 ), .B(
        \U1/aes_core/SB1/n3008 ), .C(\U1/aes_core/SB1/n3007 ), .D(
        \U1/aes_core/SB1/n3006 ), .E(\U1/aes_core/SB1/n3005 ), .F(
        \U1/aes_core/SB1/n3004 ), .Y(\U1/aes_core/SB1/n3109 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U132  ( .A0(\U1/aes_core/SB1/n3196 ), 
        .A1(\U1/aes_core/SB1/n3113 ), .B0(\U1/aes_core/SB1/n3010 ), .Y(
        \U1/aes_core/SB1/n3025 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U131  ( .AN(\U1/aes_core/SB1/n3014 ), 
        .B(\U1/aes_core/SB1/n3013 ), .C(\U1/aes_core/SB1/n3012 ), .D(
        \U1/aes_core/SB1/n3011 ), .Y(\U1/aes_core/SB1/n3024 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U130  ( .A(\U1/aes_core/SB1/n3230 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3244 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U129  ( .A(\U1/aes_core/SB1/n3017 ), .B(
        \U1/aes_core/SB1/n3016 ), .C(\U1/aes_core/SB1/n3015 ), .D(
        \U1/aes_core/SB1/n3244 ), .Y(\U1/aes_core/SB1/n3023 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U128  ( .A(\U1/aes_core/SB1/n3021 ), .B(
        \U1/aes_core/SB1/n3020 ), .C(\U1/aes_core/SB1/n3019 ), .D(
        \U1/aes_core/SB1/n3018 ), .Y(\U1/aes_core/SB1/n3022 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U127  ( .A(\U1/aes_core/SB1/n3027 ), .B(
        \U1/aes_core/SB1/n3026 ), .C(\U1/aes_core/SB1/n3025 ), .D(
        \U1/aes_core/SB1/n3024 ), .E(\U1/aes_core/SB1/n3023 ), .F(
        \U1/aes_core/SB1/n3022 ), .Y(\U1/aes_core/SB1/n3133 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U126  ( .AN(\U1/aes_core/SB1/n3031 ), 
        .B(\U1/aes_core/SB1/n3030 ), .C(\U1/aes_core/SB1/n3029 ), .D(
        \U1/aes_core/SB1/n3028 ), .Y(\U1/aes_core/SB1/n3040 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U125  ( .A(\U1/aes_core/SB1/n3035 ), .B(
        \U1/aes_core/SB1/n3034 ), .C(\U1/aes_core/SB1/n3033 ), .D(
        \U1/aes_core/SB1/n3032 ), .Y(\U1/aes_core/SB1/n3039 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U124  ( .A(\U1/aes_core/SB1/n3195 ), .B(
        \U1/aes_core/SB1/n3231 ), .C(\U1/aes_core/SB1/n3233 ), .Y(
        \U1/aes_core/SB1/n3037 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U123  ( .A0(\U1/aes_core/SB1/n3037 ), 
        .A1(\U1/aes_core/SB1/n3221 ), .B0(\U1/aes_core/SB1/n3076 ), .B1(
        \U1/aes_core/SB1/n3257 ), .C0(\U1/aes_core/SB1/n3036 ), .Y(
        \U1/aes_core/SB1/n3038 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U122  ( .A(\U1/aes_core/SB1/n3043 ), .B(
        \U1/aes_core/SB1/n3042 ), .C(\U1/aes_core/SB1/n3041 ), .D(
        \U1/aes_core/SB1/n3040 ), .E(\U1/aes_core/SB1/n3039 ), .F(
        \U1/aes_core/SB1/n3038 ), .Y(\U1/aes_core/SB1/n3181 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U121  ( .A0(\U1/aes_core/SB1/n3076 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3044 ), .Y(
        \U1/aes_core/SB1/n3058 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U120  ( .A0(\U1/aes_core/SB1/n3185 ), 
        .A1(\U1/aes_core/SB1/n3187 ), .B0(\U1/aes_core/SB1/n3242 ), .B1(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3045 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U119  ( .A0(\U1/aes_core/SB1/n3096 ), 
        .A1(\U1/aes_core/SB1/n3184 ), .B0(\U1/aes_core/SB1/n3097 ), .B1(
        \U1/aes_core/SB1/n3161 ), .C0(\U1/aes_core/SB1/n3045 ), .Y(
        \U1/aes_core/SB1/n3057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U118  ( .A(\U1/aes_core/SB1/n3046 ), .Y(
        \U1/aes_core/SB1/n3049 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U117  ( .AN(\U1/aes_core/SB1/n3050 ), 
        .B(\U1/aes_core/SB1/n3049 ), .C(\U1/aes_core/SB1/n3048 ), .D(
        \U1/aes_core/SB1/n3047 ), .Y(\U1/aes_core/SB1/n3056 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U116  ( .A(\U1/aes_core/SB1/n3054 ), .B(
        \U1/aes_core/SB1/n3053 ), .C(\U1/aes_core/SB1/n3052 ), .D(
        \U1/aes_core/SB1/n3051 ), .Y(\U1/aes_core/SB1/n3055 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U115  ( .A(\U1/aes_core/SB1/n3060 ), .B(
        \U1/aes_core/SB1/n3059 ), .C(\U1/aes_core/SB1/n3058 ), .D(
        \U1/aes_core/SB1/n3057 ), .E(\U1/aes_core/SB1/n3056 ), .F(
        \U1/aes_core/SB1/n3055 ), .Y(\U1/aes_core/SB1/n3140 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U114  ( .A0(\U1/aes_core/SB1/n3231 ), 
        .A1(\U1/aes_core/SB1/n3061 ), .B0(\U1/aes_core/SB1/n3241 ), .B1(
        \U1/aes_core/SB1/n3187 ), .Y(\U1/aes_core/SB1/n3062 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U113  ( .A0(\U1/aes_core/SB1/n3113 ), 
        .A1(\U1/aes_core/SB1/n3258 ), .B0(\U1/aes_core/SB1/n3063 ), .B1(
        \U1/aes_core/SB1/n3248 ), .C0(\U1/aes_core/SB1/n3062 ), .Y(
        \U1/aes_core/SB1/n3075 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U112  ( .AN(\U1/aes_core/SB1/n3067 ), 
        .B(\U1/aes_core/SB1/n3066 ), .C(\U1/aes_core/SB1/n3065 ), .D(
        \U1/aes_core/SB1/n3064 ), .Y(\U1/aes_core/SB1/n3074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U111  ( .A0(\U1/aes_core/SB1/n3251 ), 
        .A1(\U1/aes_core/SB1/n3068 ), .B0(\U1/aes_core/SB1/n3242 ), .Y(
        \U1/aes_core/SB1/n3072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U110  ( .A(\U1/aes_core/SB1/n3218 ), .B(
        \U1/aes_core/SB1/n3223 ), .Y(\U1/aes_core/SB1/n3069 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U109  ( .A0(\U1/aes_core/SB1/n3194 ), 
        .A1(\U1/aes_core/SB1/n3069 ), .B0(\U1/aes_core/SB1/n3195 ), .B1(
        \U1/aes_core/SB1/n3141 ), .Y(\U1/aes_core/SB1/n3070 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U108  ( .A(\U1/aes_core/SB1/n3072 ), .B(
        \U1/aes_core/SB1/n3071 ), .C(\U1/aes_core/SB1/n3070 ), .Y(
        \U1/aes_core/SB1/n3073 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U107  ( .A(\U1/aes_core/SB1/n3133 ), .B(
        \U1/aes_core/SB1/n3181 ), .C(\U1/aes_core/SB1/n3140 ), .D(
        \U1/aes_core/SB1/n3075 ), .E(\U1/aes_core/SB1/n3074 ), .F(
        \U1/aes_core/SB1/n3073 ), .Y(\U1/aes_core/SB1/n3227 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U106  ( .A(\U1/aes_core/SB1/n3160 ), .B(
        \U1/aes_core/SB1/n3205 ), .C(\U1/aes_core/SB1/n3109 ), .D(
        \U1/aes_core/SB1/n3227 ), .Y(\U1/aes_core/SB1/n3089 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U105  ( .A0(\U1/aes_core/SB1/n3207 ), 
        .A1(\U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3076 ), .B1(
        \U1/aes_core/SB1/n3223 ), .Y(\U1/aes_core/SB1/n3077 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U104  ( .A0(\U1/aes_core/SB1/n3212 ), 
        .A1(\U1/aes_core/SB1/n3230 ), .B0(\U1/aes_core/SB1/n3243 ), .B1(
        \U1/aes_core/SB1/n3251 ), .C0(\U1/aes_core/SB1/n3077 ), .Y(
        \U1/aes_core/SB1/n3088 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U103  ( .A(\U1/aes_core/SB1/n3078 ), .Y(
        \U1/aes_core/SB1/n3081 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U102  ( .A0(\U1/aes_core/SB1/n3079 ), 
        .A1(\U1/aes_core/SB1/n3184 ), .B0(\U1/aes_core/SB1/n3112 ), .B1(
        \U1/aes_core/SB1/n3164 ), .Y(\U1/aes_core/SB1/n3080 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U101  ( .A0(\U1/aes_core/SB1/n3231 ), 
        .A1(\U1/aes_core/SB1/n3081 ), .B0(\U1/aes_core/SB1/n3213 ), .B1(
        \U1/aes_core/SB1/n3162 ), .C0(\U1/aes_core/SB1/n3080 ), .Y(
        \U1/aes_core/SB1/n3087 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U100  ( .A0(\U1/aes_core/SB1/n3253 ), 
        .A1(\U1/aes_core/SB1/n3130 ), .B0(\U1/aes_core/SB1/n3233 ), .Y(
        \U1/aes_core/SB1/n3085 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB1/U99  ( .A(\U1/aes_core/SB1/n3085 ), .B(
        \U1/aes_core/SB1/n3084 ), .C(\U1/aes_core/SB1/n3083 ), .D(
        \U1/aes_core/SB1/n3082 ), .Y(\U1/aes_core/SB1/n3086 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U98  ( .AN(\U1/aes_core/SB1/n3089 ), .B(
        \U1/aes_core/SB1/n3088 ), .C(\U1/aes_core/SB1/n3087 ), .D(
        \U1/aes_core/SB1/n3086 ), .Y(\U1/aes_core/sb1 [3]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U97  ( .A0(\U1/aes_core/SB1/n3104 ), .A1(
        \U1/aes_core/SB1/n3219 ), .B0(\U1/aes_core/SB1/n3163 ), .Y(
        \U1/aes_core/SB1/n3101 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U96  ( .A(\U1/aes_core/SB1/n3092 ), .B(
        \U1/aes_core/SB1/n3091 ), .C(\U1/aes_core/SB1/n3090 ), .Y(
        \U1/aes_core/SB1/n3100 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U95  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3242 ), .Y(\U1/aes_core/SB1/n3095 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U94  ( .A(\U1/aes_core/SB1/n3213 ), .B(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3093 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U93  ( .A0(\U1/aes_core/SB1/n3095 ), 
        .A1(\U1/aes_core/SB1/n3094 ), .B0(\U1/aes_core/SB1/n3093 ), .B1(
        \U1/aes_core/SB1/n3236 ), .C0(\U1/aes_core/SB1/n3219 ), .C1(
        \U1/aes_core/SB1/n3145 ), .Y(\U1/aes_core/SB1/n3099 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U92  ( .A0(\U1/aes_core/SB1/n3196 ), 
        .A1(\U1/aes_core/SB1/n3097 ), .B0(\U1/aes_core/SB1/n3258 ), .B1(
        \U1/aes_core/SB1/n3248 ), .C0(\U1/aes_core/SB1/n3221 ), .C1(
        \U1/aes_core/SB1/n3096 ), .Y(\U1/aes_core/SB1/n3098 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U91  ( .A(\U1/aes_core/SB1/n3103 ), .B(
        \U1/aes_core/SB1/n3102 ), .C(\U1/aes_core/SB1/n3101 ), .D(
        \U1/aes_core/SB1/n3100 ), .E(\U1/aes_core/SB1/n3099 ), .F(
        \U1/aes_core/SB1/n3098 ), .Y(\U1/aes_core/SB1/n3228 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB1/U90  ( .A0(\U1/aes_core/SB1/n3104 ), .A1(
        \U1/aes_core/SB1/n3113 ), .B0(\U1/aes_core/SB1/n3184 ), .Y(
        \U1/aes_core/SB1/n3139 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB1/U89  ( .A0(\U1/aes_core/SB1/n3208 ), .A1(
        \U1/aes_core/SB1/n3221 ), .A2(\U1/aes_core/SB1/n3161 ), .B0(
        \U1/aes_core/SB1/n3237 ), .Y(\U1/aes_core/SB1/n3138 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U88  ( .A(\U1/aes_core/SB1/n3108 ), .B(
        \U1/aes_core/SB1/n3107 ), .C(\U1/aes_core/SB1/n3106 ), .D(
        \U1/aes_core/SB1/n3105 ), .Y(\U1/aes_core/SB1/n3135 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U87  ( .A(\U1/aes_core/SB1/n3109 ), .Y(
        \U1/aes_core/SB1/n3132 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U86  ( .A(\U1/aes_core/SB1/n3110 ), .Y(
        \U1/aes_core/SB1/n3126 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB1/U85  ( .A0(\U1/aes_core/SB1/n3112 ), 
        .A1(\U1/aes_core/SB1/n3249 ), .B0N(\U1/aes_core/SB1/n3111 ), .Y(
        \U1/aes_core/SB1/n3125 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U84  ( .A0(\U1/aes_core/SB1/n3256 ), 
        .A1(\U1/aes_core/SB1/n3113 ), .B0(\U1/aes_core/SB1/n3163 ), .B1(
        \U1/aes_core/SB1/n3223 ), .C0(\U1/aes_core/SB1/n3237 ), .C1(
        \U1/aes_core/SB1/n3258 ), .Y(\U1/aes_core/SB1/n3124 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U83  ( .AN(\U1/aes_core/SB1/n3117 ), .B(
        \U1/aes_core/SB1/n3116 ), .C(\U1/aes_core/SB1/n3115 ), .D(
        \U1/aes_core/SB1/n3114 ), .Y(\U1/aes_core/SB1/n3123 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U82  ( .A(\U1/aes_core/SB1/n3121 ), .B(
        \U1/aes_core/SB1/n3120 ), .C(\U1/aes_core/SB1/n3119 ), .D(
        \U1/aes_core/SB1/n3118 ), .Y(\U1/aes_core/SB1/n3122 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U81  ( .A(\U1/aes_core/SB1/n3127 ), .B(
        \U1/aes_core/SB1/n3126 ), .C(\U1/aes_core/SB1/n3125 ), .D(
        \U1/aes_core/SB1/n3124 ), .E(\U1/aes_core/SB1/n3123 ), .F(
        \U1/aes_core/SB1/n3122 ), .Y(\U1/aes_core/SB1/n3128 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U80  ( .A(\U1/aes_core/SB1/n3128 ), .Y(
        \U1/aes_core/SB1/n3206 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U79  ( .A0(\U1/aes_core/SB1/n3196 ), .A1(
        \U1/aes_core/SB1/n3218 ), .B0(\U1/aes_core/SB1/n3258 ), .B1(
        \U1/aes_core/SB1/n3257 ), .Y(\U1/aes_core/SB1/n3129 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U78  ( .A0(\U1/aes_core/SB1/n3186 ), 
        .A1(\U1/aes_core/SB1/n3130 ), .B0(\U1/aes_core/SB1/n3210 ), .B1(
        \U1/aes_core/SB1/n3232 ), .C0(\U1/aes_core/SB1/n3129 ), .Y(
        \U1/aes_core/SB1/n3131 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U77  ( .AN(\U1/aes_core/SB1/n3133 ), .B(
        \U1/aes_core/SB1/n3132 ), .C(\U1/aes_core/SB1/n3206 ), .D(
        \U1/aes_core/SB1/n3131 ), .Y(\U1/aes_core/SB1/n3134 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U76  ( .A(\U1/aes_core/SB1/n3139 ), .B(
        \U1/aes_core/SB1/n3138 ), .C(\U1/aes_core/SB1/n3137 ), .D(
        \U1/aes_core/SB1/n3136 ), .E(\U1/aes_core/SB1/n3135 ), .F(
        \U1/aes_core/SB1/n3134 ), .Y(\U1/aes_core/SB1/n3204 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U75  ( .A(\U1/aes_core/SB1/n3140 ), .Y(
        \U1/aes_core/SB1/n3144 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U74  ( .A0(\U1/aes_core/SB1/n3142 ), .A1(
        \U1/aes_core/SB1/n3141 ), .B0(\U1/aes_core/SB1/n3188 ), .B1(
        \U1/aes_core/SB1/n3147 ), .Y(\U1/aes_core/SB1/n3143 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U73  ( .A0(\U1/aes_core/SB1/n3237 ), 
        .A1(\U1/aes_core/SB1/n3145 ), .B0(\U1/aes_core/SB1/n3144 ), .C0(
        \U1/aes_core/SB1/n3143 ), .Y(\U1/aes_core/SB1/n3159 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U72  ( .A0(\U1/aes_core/SB1/n3146 ), .A1(
        \U1/aes_core/SB1/n3209 ), .B0(\U1/aes_core/SB1/n3238 ), .Y(
        \U1/aes_core/SB1/n3151 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U71  ( .A0(\U1/aes_core/SB1/n3147 ), .A1(
        \U1/aes_core/SB1/n3212 ), .B0(\U1/aes_core/SB1/n3241 ), .Y(
        \U1/aes_core/SB1/n3150 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U70  ( .A(\U1/aes_core/SB1/n3151 ), .B(
        \U1/aes_core/SB1/n3150 ), .C(\U1/aes_core/SB1/n3149 ), .D(
        \U1/aes_core/SB1/n3148 ), .Y(\U1/aes_core/SB1/n3158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U69  ( .A(\U1/aes_core/SB1/n3189 ), .B(
        \U1/aes_core/SB1/n3152 ), .Y(\U1/aes_core/SB1/n3156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U68  ( .A(\U1/aes_core/SB1/n3153 ), .B(
        \U1/aes_core/SB1/n3194 ), .Y(\U1/aes_core/SB1/n3155 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U67  ( .A0(\U1/aes_core/SB1/n3156 ), 
        .A1(\U1/aes_core/SB1/n3255 ), .B0(\U1/aes_core/SB1/n3155 ), .B1(
        \U1/aes_core/SB1/n3219 ), .C0(\U1/aes_core/SB1/n3154 ), .C1(
        \U1/aes_core/SB1/n3220 ), .Y(\U1/aes_core/SB1/n3157 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U66  ( .A(\U1/aes_core/SB1/n3228 ), .B(
        \U1/aes_core/SB1/n3204 ), .C(\U1/aes_core/SB1/n3160 ), .D(
        \U1/aes_core/SB1/n3159 ), .E(\U1/aes_core/SB1/n3158 ), .F(
        \U1/aes_core/SB1/n3157 ), .Y(\U1/aes_core/sb1 [4]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U65  ( .A1N(\U1/aes_core/SB1/n3162 ), 
        .A0(\U1/aes_core/SB1/n3161 ), .B0(\U1/aes_core/SB1/n3218 ), .Y(
        \U1/aes_core/SB1/n3178 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U64  ( .A(\U1/aes_core/SB1/n3231 ), .B(
        \U1/aes_core/SB1/n3212 ), .Y(\U1/aes_core/SB1/n3165 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U63  ( .A0(\U1/aes_core/SB1/n3255 ), 
        .A1(\U1/aes_core/SB1/n3166 ), .B0(\U1/aes_core/SB1/n3165 ), .B1(
        \U1/aes_core/SB1/n3258 ), .C0(\U1/aes_core/SB1/n3164 ), .C1(
        \U1/aes_core/SB1/n3163 ), .Y(\U1/aes_core/SB1/n3177 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U62  ( .A(\U1/aes_core/SB1/n3167 ), .Y(
        \U1/aes_core/SB1/n3170 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U61  ( .AN(\U1/aes_core/SB1/n3171 ), .B(
        \U1/aes_core/SB1/n3170 ), .C(\U1/aes_core/SB1/n3169 ), .D(
        \U1/aes_core/SB1/n3168 ), .Y(\U1/aes_core/SB1/n3176 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U60  ( .A(\U1/aes_core/SB1/n3174 ), .B(
        \U1/aes_core/SB1/n3173 ), .C(\U1/aes_core/SB1/n3172 ), .Y(
        \U1/aes_core/SB1/n3175 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U59  ( .A(\U1/aes_core/SB1/n3180 ), .B(
        \U1/aes_core/SB1/n3179 ), .C(\U1/aes_core/SB1/n3178 ), .D(
        \U1/aes_core/SB1/n3177 ), .E(\U1/aes_core/SB1/n3176 ), .F(
        \U1/aes_core/SB1/n3175 ), .Y(\U1/aes_core/SB1/n3229 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U58  ( .A(\U1/aes_core/SB1/n3181 ), .Y(
        \U1/aes_core/SB1/n3183 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U57  ( .A0(\U1/aes_core/SB1/n3242 ), .A1(
        \U1/aes_core/SB1/n3239 ), .B0(\U1/aes_core/SB1/n3243 ), .B1(
        \U1/aes_core/SB1/n3241 ), .Y(\U1/aes_core/SB1/n3182 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U56  ( .A0(\U1/aes_core/SB1/n3218 ), 
        .A1(\U1/aes_core/SB1/n3184 ), .B0(\U1/aes_core/SB1/n3183 ), .C0(
        \U1/aes_core/SB1/n3182 ), .Y(\U1/aes_core/SB1/n3203 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U55  ( .A0(\U1/aes_core/SB1/n3186 ), .A1(
        \U1/aes_core/SB1/n3242 ), .B0(\U1/aes_core/SB1/n3185 ), .Y(
        \U1/aes_core/SB1/n3192 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U54  ( .A0(\U1/aes_core/SB1/n3189 ), .A1(
        \U1/aes_core/SB1/n3188 ), .B0(\U1/aes_core/SB1/n3187 ), .Y(
        \U1/aes_core/SB1/n3191 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U53  ( .AN(\U1/aes_core/SB1/n3193 ), .B(
        \U1/aes_core/SB1/n3192 ), .C(\U1/aes_core/SB1/n3191 ), .D(
        \U1/aes_core/SB1/n3190 ), .Y(\U1/aes_core/SB1/n3202 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U52  ( .A0(\U1/aes_core/SB1/n3238 ), .A1(
        \U1/aes_core/SB1/n3195 ), .B0(\U1/aes_core/SB1/n3194 ), .Y(
        \U1/aes_core/SB1/n3199 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB1/U51  ( .A0(\U1/aes_core/SB1/n3220 ), .A1(
        \U1/aes_core/SB1/n3197 ), .B0(\U1/aes_core/SB1/n3257 ), .B1(
        \U1/aes_core/SB1/n3196 ), .Y(\U1/aes_core/SB1/n3198 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U50  ( .A0(\U1/aes_core/SB1/n3200 ), 
        .A1(\U1/aes_core/SB1/n3219 ), .B0(\U1/aes_core/SB1/n3199 ), .C0(
        \U1/aes_core/SB1/n3198 ), .Y(\U1/aes_core/SB1/n3201 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U49  ( .A(\U1/aes_core/SB1/n3229 ), .B(
        \U1/aes_core/SB1/n3205 ), .C(\U1/aes_core/SB1/n3204 ), .D(
        \U1/aes_core/SB1/n3203 ), .E(\U1/aes_core/SB1/n3202 ), .F(
        \U1/aes_core/SB1/n3201 ), .Y(\U1/aes_core/sb1 [5]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U48  ( .A0(\U1/aes_core/SB1/n3208 ), 
        .A1(\U1/aes_core/SB1/n3248 ), .B0(\U1/aes_core/SB1/n3207 ), .B1(
        \U1/aes_core/SB1/n3255 ), .C0(\U1/aes_core/SB1/n3206 ), .Y(
        \U1/aes_core/SB1/n3226 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U47  ( .A0(\U1/aes_core/SB1/n3209 ), .A1(
        \U1/aes_core/SB1/n3253 ), .B0(\U1/aes_core/SB1/n3242 ), .Y(
        \U1/aes_core/SB1/n3217 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U46  ( .A0(\U1/aes_core/SB1/n3233 ), .A1(
        \U1/aes_core/SB1/n3210 ), .B0(\U1/aes_core/SB1/n3241 ), .Y(
        \U1/aes_core/SB1/n3216 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U45  ( .A0(\U1/aes_core/SB1/n3213 ), .A1(
        \U1/aes_core/SB1/n3212 ), .B0(\U1/aes_core/SB1/n3211 ), .Y(
        \U1/aes_core/SB1/n3215 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U44  ( .A(\U1/aes_core/SB1/n3217 ), .B(
        \U1/aes_core/SB1/n3216 ), .C(\U1/aes_core/SB1/n3215 ), .D(
        \U1/aes_core/SB1/n3214 ), .Y(\U1/aes_core/SB1/n3225 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U43  ( .A(\U1/aes_core/SB1/n3248 ), .B(
        \U1/aes_core/SB1/n3218 ), .Y(\U1/aes_core/SB1/n3250 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB1/U42  ( .A(\U1/aes_core/SB1/n3238 ), .B(
        \U1/aes_core/SB1/n3250 ), .Y(\U1/aes_core/SB1/n3222 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U41  ( .A0(\U1/aes_core/SB1/n3236 ), 
        .A1(\U1/aes_core/SB1/n3223 ), .B0(\U1/aes_core/SB1/n3222 ), .B1(
        \U1/aes_core/SB1/n3221 ), .C0(\U1/aes_core/SB1/n3220 ), .C1(
        \U1/aes_core/SB1/n3219 ), .Y(\U1/aes_core/SB1/n3224 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U40  ( .A(\U1/aes_core/SB1/n3229 ), .B(
        \U1/aes_core/SB1/n3228 ), .C(\U1/aes_core/SB1/n3227 ), .D(
        \U1/aes_core/SB1/n3226 ), .E(\U1/aes_core/SB1/n3225 ), .F(
        \U1/aes_core/SB1/n3224 ), .Y(\U1/aes_core/sb1 [6]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U39  ( .A0(\U1/aes_core/SB1/n3233 ), .A1(
        \U1/aes_core/SB1/n3232 ), .B0(\U1/aes_core/SB1/n3231 ), .B1(
        \U1/aes_core/SB1/n3230 ), .Y(\U1/aes_core/SB1/n3234 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB1/U38  ( .A0(\U1/aes_core/SB1/n3237 ), 
        .A1(\U1/aes_core/SB1/n3236 ), .B0(\U1/aes_core/SB1/n3235 ), .C0(
        \U1/aes_core/SB1/n3234 ), .Y(\U1/aes_core/SB1/n3261 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB1/U37  ( .A1N(\U1/aes_core/SB1/n3240 ), 
        .A0(\U1/aes_core/SB1/n3239 ), .B0(\U1/aes_core/SB1/n3238 ), .Y(
        \U1/aes_core/SB1/n3247 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U36  ( .A0(\U1/aes_core/SB1/n3243 ), .A1(
        \U1/aes_core/SB1/n3242 ), .B0(\U1/aes_core/SB1/n3241 ), .Y(
        \U1/aes_core/SB1/n3246 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U35  ( .A(\U1/aes_core/SB1/n3247 ), .B(
        \U1/aes_core/SB1/n3246 ), .C(\U1/aes_core/SB1/n3245 ), .D(
        \U1/aes_core/SB1/n3244 ), .Y(\U1/aes_core/SB1/n3260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U34  ( .A(\U1/aes_core/SB1/n3249 ), .B(
        \U1/aes_core/SB1/n3248 ), .Y(\U1/aes_core/SB1/n3252 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U33  ( .A0(\U1/aes_core/SB1/n3253 ), .A1(
        \U1/aes_core/SB1/n3252 ), .B0(\U1/aes_core/SB1/n3251 ), .B1(
        \U1/aes_core/SB1/n3250 ), .Y(\U1/aes_core/SB1/n3254 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U32  ( .A0(\U1/aes_core/SB1/n3258 ), 
        .A1(\U1/aes_core/SB1/n3257 ), .B0(\U1/aes_core/SB1/n3256 ), .B1(
        \U1/aes_core/SB1/n3255 ), .C0(\U1/aes_core/SB1/n3254 ), .Y(
        \U1/aes_core/SB1/n3259 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U31  ( .A(\U1/aes_core/SB1/n3264 ), .B(
        \U1/aes_core/SB1/n3263 ), .C(\U1/aes_core/SB1/n3262 ), .D(
        \U1/aes_core/SB1/n3261 ), .E(\U1/aes_core/SB1/n3260 ), .F(
        \U1/aes_core/SB1/n3259 ), .Y(\U1/aes_core/sb1 [7]) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U30  ( .A(\U1/aes_core/SB1/n3267 ), .B(
        \U1/aes_core/SB1/n3266 ), .C(\U1/aes_core/SB1/n3265 ), .Y(
        \U1/aes_core/SB1/n3290 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U29  ( .A0(\U1/aes_core/SB1/n3268 ), .A1(
        \U1/aes_core/SB1/n3324 ), .B0(\U1/aes_core/SB1/n3340 ), .Y(
        \U1/aes_core/SB1/n3273 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U28  ( .A0(\U1/aes_core/SB1/n3333 ), .A1(
        \U1/aes_core/SB1/n3270 ), .B0(\U1/aes_core/SB1/n3269 ), .B1(
        \U1/aes_core/SB1/n3334 ), .Y(\U1/aes_core/SB1/n3271 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U27  ( .A(\U1/aes_core/SB1/n3273 ), .B(
        \U1/aes_core/SB1/n3272 ), .C(\U1/aes_core/SB1/n3271 ), .Y(
        \U1/aes_core/SB1/n3289 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB1/U26  ( .A0(\U1/aes_core/SB1/n3276 ), .A1(
        \U1/aes_core/SB1/n3299 ), .B0(\U1/aes_core/SB1/n3275 ), .B1(
        \U1/aes_core/SB1/n3274 ), .Y(\U1/aes_core/SB1/n3277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB1/U25  ( .A0(\U1/aes_core/SB1/n3281 ), 
        .A1(\U1/aes_core/SB1/n3280 ), .B0(\U1/aes_core/SB1/n3279 ), .B1(
        \U1/aes_core/SB1/n3278 ), .C0(\U1/aes_core/SB1/n3277 ), .Y(
        \U1/aes_core/SB1/n3288 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U24  ( .A(\U1/aes_core/SB1/n3329 ), .B(
        \U1/aes_core/SB1/n3282 ), .Y(\U1/aes_core/SB1/n3283 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U23  ( .AN(\U1/aes_core/SB1/n3286 ), .B(
        \U1/aes_core/SB1/n3285 ), .C(\U1/aes_core/SB1/n3284 ), .D(
        \U1/aes_core/SB1/n3283 ), .Y(\U1/aes_core/SB1/n3287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U22  ( .A(\U1/aes_core/SB1/n3292 ), .B(
        \U1/aes_core/SB1/n3291 ), .C(\U1/aes_core/SB1/n3290 ), .D(
        \U1/aes_core/SB1/n3289 ), .E(\U1/aes_core/SB1/n3288 ), .F(
        \U1/aes_core/SB1/n3287 ), .Y(\U1/aes_core/SB1/n3351 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB1/U21  ( .A(\U1/aes_core/SB1/n3295 ), .B(
        \U1/aes_core/SB1/n3294 ), .C(\U1/aes_core/SB1/n3293 ), .D(
        \U1/aes_core/SB1/n3351 ), .Y(\U1/aes_core/SB1/n3320 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U20  ( .A0(\U1/aes_core/SB1/n3297 ), .A1(
        \U1/aes_core/SB1/n3308 ), .B0(\U1/aes_core/SB1/n3344 ), .B1(
        \U1/aes_core/SB1/n3296 ), .Y(\U1/aes_core/SB1/n3298 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U19  ( .A0(\U1/aes_core/SB1/n3322 ), 
        .A1(\U1/aes_core/SB1/n3334 ), .B0(\U1/aes_core/SB1/n3325 ), .B1(
        \U1/aes_core/SB1/n3299 ), .C0(\U1/aes_core/SB1/n3298 ), .Y(
        \U1/aes_core/SB1/n3319 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB1/U18  ( .A0(\U1/aes_core/SB1/n3303 ), .A1(
        \U1/aes_core/SB1/n3302 ), .B0(\U1/aes_core/SB1/n3301 ), .B1(
        \U1/aes_core/SB1/n3300 ), .Y(\U1/aes_core/SB1/n3304 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U17  ( .A0(\U1/aes_core/SB1/n3307 ), 
        .A1(\U1/aes_core/SB1/n3306 ), .B0(\U1/aes_core/SB1/n3305 ), .B1(
        \U1/aes_core/SB1/n3330 ), .C0(\U1/aes_core/SB1/n3304 ), .Y(
        \U1/aes_core/SB1/n3318 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB1/U16  ( .A(\U1/aes_core/SB1/n3309 ), .B(
        \U1/aes_core/SB1/n3308 ), .Y(\U1/aes_core/SB1/n3316 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U15  ( .A(\U1/aes_core/SB1/n3310 ), .Y(
        \U1/aes_core/SB1/n3315 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB1/U14  ( .A(\U1/aes_core/SB1/n3313 ), .B(
        \U1/aes_core/SB1/n3312 ), .C(\U1/aes_core/SB1/n3311 ), .Y(
        \U1/aes_core/SB1/n3314 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U13  ( .A0(\U1/aes_core/SB1/n3331 ), 
        .A1(\U1/aes_core/SB1/n3316 ), .B0(\U1/aes_core/SB1/n3323 ), .B1(
        \U1/aes_core/SB1/n3315 ), .C0(\U1/aes_core/SB1/n3314 ), .Y(
        \U1/aes_core/SB1/n3317 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB1/U12  ( .AN(\U1/aes_core/SB1/n3320 ), .B(
        \U1/aes_core/SB1/n3319 ), .C(\U1/aes_core/SB1/n3318 ), .D(
        \U1/aes_core/SB1/n3317 ), .Y(\U1/aes_core/sb1 [8]) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB1/U11  ( .A0(\U1/aes_core/SB1/n3325 ), 
        .A1(\U1/aes_core/SB1/n3324 ), .B0(\U1/aes_core/SB1/n3323 ), .B1(
        \U1/aes_core/SB1/n3322 ), .C0(\U1/aes_core/SB1/n3321 ), .Y(
        \U1/aes_core/SB1/n3326 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB1/U10  ( .A(\U1/aes_core/SB1/n3326 ), .Y(
        \U1/aes_core/SB1/n3350 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U9  ( .A0(\U1/aes_core/SB1/n3339 ), .A1(
        \U1/aes_core/SB1/n3328 ), .B0(\U1/aes_core/SB1/n3327 ), .Y(
        \U1/aes_core/SB1/n3338 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U8  ( .A0(\U1/aes_core/SB1/n3331 ), .A1(
        \U1/aes_core/SB1/n3330 ), .B0(\U1/aes_core/SB1/n3329 ), .Y(
        \U1/aes_core/SB1/n3337 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB1/U7  ( .A0(\U1/aes_core/SB1/n3334 ), .A1(
        \U1/aes_core/SB1/n3333 ), .B0(\U1/aes_core/SB1/n3332 ), .Y(
        \U1/aes_core/SB1/n3336 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB1/U6  ( .A(\U1/aes_core/SB1/n3338 ), .B(
        \U1/aes_core/SB1/n3337 ), .C(\U1/aes_core/SB1/n3336 ), .D(
        \U1/aes_core/SB1/n3335 ), .Y(\U1/aes_core/SB1/n3349 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB1/U5  ( .A(\U1/aes_core/SB1/n3341 ), .B(
        \U1/aes_core/SB1/n3340 ), .C(\U1/aes_core/SB1/n3339 ), .Y(
        \U1/aes_core/SB1/n3345 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB1/U4  ( .A0(\U1/aes_core/SB1/n3347 ), .A1(
        \U1/aes_core/SB1/n3346 ), .B0(\U1/aes_core/SB1/n3345 ), .B1(
        \U1/aes_core/SB1/n3344 ), .C0(\U1/aes_core/SB1/n3343 ), .C1(
        \U1/aes_core/SB1/n3342 ), .Y(\U1/aes_core/SB1/n3348 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB1/U3  ( .A(\U1/aes_core/SB1/n3353 ), .B(
        \U1/aes_core/SB1/n3352 ), .C(\U1/aes_core/SB1/n3351 ), .D(
        \U1/aes_core/SB1/n3350 ), .E(\U1/aes_core/SB1/n3349 ), .F(
        \U1/aes_core/SB1/n3348 ), .Y(\U1/aes_core/sb1 [9]) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U711  ( .A0(\U1/aes_core/SB2/n2203 ), .A1(
        \U1/aes_core/SB2/n2353 ), .B0(\U1/aes_core/SB2/n2351 ), .B1(
        \U1/aes_core/SB2/n2311 ), .C0(\U1/aes_core/SB2/n2202 ), .Y(
        \U1/aes_core/SB2/n2205 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U393  ( .A0(\U1/aes_core/SB2/n2650 ), .A1(
        \U1/aes_core/SB2/n2775 ), .B0(\U1/aes_core/SB2/n2773 ), .B1(
        \U1/aes_core/SB2/n2758 ), .C0(\U1/aes_core/SB2/n2649 ), .Y(
        \U1/aes_core/SB2/n2652 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U391  ( .A0(\U1/aes_core/SB2/n3145 ), .A1(
        \U1/aes_core/SB2/n2328 ), .B0(\U1/aes_core/SB2/n3223 ), .B1(
        \U1/aes_core/SB2/n3207 ), .C0(\U1/aes_core/SB2/n2993 ), .Y(
        \U1/aes_core/SB2/n2329 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U363  ( .A0(\U1/aes_core/SB2/n2402 ), .A1(
        \U1/aes_core/SB2/n2157 ), .B0(\U1/aes_core/SB2/n2480 ), .B1(
        \U1/aes_core/SB2/n2464 ), .C0(\U1/aes_core/SB2/n2225 ), .Y(
        \U1/aes_core/SB2/n2158 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U361  ( .A0(\U1/aes_core/SB2/n2824 ), .A1(
        \U1/aes_core/SB2/n2604 ), .B0(\U1/aes_core/SB2/n2923 ), .B1(
        \U1/aes_core/SB2/n2907 ), .C0(\U1/aes_core/SB2/n2672 ), .Y(
        \U1/aes_core/SB2/n2605 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U301  ( .A0(\U1/aes_core/SB2/n2971 ), .A1(
        \U1/aes_core/SB2/n3096 ), .B0(\U1/aes_core/SB2/n3094 ), .B1(
        \U1/aes_core/SB2/n3079 ), .C0(\U1/aes_core/SB2/n2970 ), .Y(
        \U1/aes_core/SB2/n2973 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U300  ( .A0(\U1/aes_core/SB2/n2402 ), .A1(
        \U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2480 ), .B1(
        \U1/aes_core/SB2/n2478 ), .C0(\U1/aes_core/SB2/n2268 ), .Y(
        \U1/aes_core/SB2/n2144 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U151  ( .A0(\U1/aes_core/SB2/n2824 ), .A1(
        \U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2923 ), .B1(
        \U1/aes_core/SB2/n2921 ), .C0(\U1/aes_core/SB2/n2715 ), .Y(
        \U1/aes_core/SB2/n2591 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB2/U150  ( .A0(\U1/aes_core/SB2/n3145 ), .A1(
        \U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3223 ), .B1(
        \U1/aes_core/SB2/n3221 ), .C0(\U1/aes_core/SB2/n3036 ), .Y(
        \U1/aes_core/SB2/n1742 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1724  ( .A(Dout[39]), .B(Dout[38]), .Y(
        \U1/aes_core/SB2/n1691 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1723  ( .A(Dout[37]), .B(Dout[36]), .Y(
        \U1/aes_core/SB2/n1682 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1722  ( .A(\U1/aes_core/SB2/n1691 ), .B(
        \U1/aes_core/SB2/n1682 ), .Y(\U1/aes_core/SB2/n2328 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1721  ( .A(Dout[33]), .Y(
        \U1/aes_core/SB2/n767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1720  ( .A(Dout[32]), .Y(
        \U1/aes_core/SB2/n385 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1719  ( .A(\U1/aes_core/SB2/n767 ), .B(
        \U1/aes_core/SB2/n385 ), .Y(\U1/aes_core/SB2/n1683 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1718  ( .A(Dout[35]), .B(Dout[34]), .Y(
        \U1/aes_core/SB2/n1703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1717  ( .A(\U1/aes_core/SB2/n1683 ), .B(
        \U1/aes_core/SB2/n1703 ), .Y(\U1/aes_core/SB2/n3207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1716  ( .A(\U1/aes_core/SB2/n2328 ), .B(
        \U1/aes_core/SB2/n3207 ), .Y(\U1/aes_core/SB2/n3014 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U1715  ( .A(Dout[34]), .B(Dout[35]), .Y(
        \U1/aes_core/SB2/n1686 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1714  ( .A(\U1/aes_core/SB2/n1686 ), .B(
        \U1/aes_core/SB2/n1683 ), .Y(\U1/aes_core/SB2/n3145 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1713  ( .A(Dout[39]), .Y(
        \U1/aes_core/SB2/n1203 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1712  ( .A(\U1/aes_core/SB2/n1203 ), .B(
        Dout[38]), .Y(\U1/aes_core/SB2/n1709 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1711  ( .A(\U1/aes_core/SB2/n1709 ), .B(
        \U1/aes_core/SB2/n1682 ), .Y(\U1/aes_core/SB2/n2327 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1710  ( .A(\U1/aes_core/SB2/n3145 ), .B(
        \U1/aes_core/SB2/n2327 ), .Y(\U1/aes_core/SB2/n3111 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1709  ( .A(Dout[35]), .Y(
        \U1/aes_core/SB2/n707 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U1708  ( .A(Dout[34]), .B(
        \U1/aes_core/SB2/n707 ), .Y(\U1/aes_core/SB2/n1684 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1707  ( .A(\U1/aes_core/SB2/n1683 ), .B(
        \U1/aes_core/SB2/n1684 ), .Y(\U1/aes_core/SB2/n3076 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1706  ( .A(\U1/aes_core/SB2/n3076 ), .Y(
        \U1/aes_core/SB2/n3241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1705  ( .A(Dout[36]), .Y(
        \U1/aes_core/SB2/n752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1704  ( .A(\U1/aes_core/SB2/n752 ), .B(
        Dout[37]), .Y(\U1/aes_core/SB2/n1690 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1703  ( .A(Dout[38]), .Y(
        \U1/aes_core/SB2/n1158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1702  ( .A(\U1/aes_core/SB2/n1158 ), .B(
        Dout[39]), .Y(\U1/aes_core/SB2/n1700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1701  ( .A(\U1/aes_core/SB2/n1690 ), .B(
        \U1/aes_core/SB2/n1700 ), .Y(\U1/aes_core/SB2/n3097 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1700  ( .A(\U1/aes_core/SB2/n3097 ), .Y(
        \U1/aes_core/SB2/n3195 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1699  ( .A(\U1/aes_core/SB2/n3241 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n3054 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1698  ( .A(\U1/aes_core/SB2/n2328 ), .Y(
        \U1/aes_core/SB2/n3210 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1697  ( .A(Dout[33]), .B(Dout[32]), .Y(
        \U1/aes_core/SB2/n1687 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1696  ( .A(\U1/aes_core/SB2/n1687 ), .B(
        \U1/aes_core/SB2/n1703 ), .Y(\U1/aes_core/SB2/n3163 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1695  ( .A(\U1/aes_core/SB2/n3163 ), .Y(
        \U1/aes_core/SB2/n3251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1694  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3251 ), .Y(\U1/aes_core/SB2/n3168 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1693  ( .A(\U1/aes_core/SB2/n385 ), .B(
        Dout[33]), .Y(\U1/aes_core/SB2/n1702 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1692  ( .A(\U1/aes_core/SB2/n1684 ), .B(
        \U1/aes_core/SB2/n1702 ), .Y(\U1/aes_core/SB2/n3063 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1691  ( .A(\U1/aes_core/SB2/n3063 ), .Y(
        \U1/aes_core/SB2/n3152 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1690  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3032 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U1689  ( .A(\U1/aes_core/SB2/n3054 ), .B(
        \U1/aes_core/SB2/n3168 ), .C(\U1/aes_core/SB2/n3032 ), .Y(
        \U1/aes_core/SB2/n1722 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1688  ( .A(\U1/aes_core/SB2/n1682 ), .B(
        \U1/aes_core/SB2/n1700 ), .Y(\U1/aes_core/SB2/n3096 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1687  ( .A(\U1/aes_core/SB2/n707 ), .B(
        Dout[34]), .Y(\U1/aes_core/SB2/n1693 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1686  ( .A(\U1/aes_core/SB2/n1693 ), .B(
        \U1/aes_core/SB2/n1702 ), .Y(\U1/aes_core/SB2/n3094 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1685  ( .A(\U1/aes_core/SB2/n3096 ), .B(
        \U1/aes_core/SB2/n3094 ), .Y(\U1/aes_core/SB2/n3009 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1684  ( .A(\U1/aes_core/SB2/n2327 ), .Y(
        \U1/aes_core/SB2/n3212 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1683  ( .A(Dout[37]), .Y(
        \U1/aes_core/SB2/n1030 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1682  ( .A(\U1/aes_core/SB2/n752 ), .B(
        \U1/aes_core/SB2/n1030 ), .Y(\U1/aes_core/SB2/n1701 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1681  ( .A(\U1/aes_core/SB2/n1691 ), .B(
        \U1/aes_core/SB2/n1701 ), .Y(\U1/aes_core/SB2/n3255 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1680  ( .A(\U1/aes_core/SB2/n3255 ), .Y(
        \U1/aes_core/SB2/n3186 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1679  ( .A(\U1/aes_core/SB2/n767 ), .B(
        Dout[32]), .Y(\U1/aes_core/SB2/n1692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1678  ( .A(\U1/aes_core/SB2/n1692 ), .B(
        \U1/aes_core/SB2/n1703 ), .Y(\U1/aes_core/SB2/n3220 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1677  ( .A(\U1/aes_core/SB2/n3220 ), .Y(
        \U1/aes_core/SB2/n3068 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1676  ( .A0(\U1/aes_core/SB2/n3212 ), 
        .A1(\U1/aes_core/SB2/n3186 ), .B0(\U1/aes_core/SB2/n3068 ), .Y(
        \U1/aes_core/SB2/n1621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1675  ( .A(\U1/aes_core/SB2/n1687 ), .B(
        \U1/aes_core/SB2/n1684 ), .Y(\U1/aes_core/SB2/n3208 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1674  ( .A(\U1/aes_core/SB2/n3208 ), .Y(
        \U1/aes_core/SB2/n3194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1673  ( .A(\U1/aes_core/SB2/n1030 ), .B(
        Dout[36]), .Y(\U1/aes_core/SB2/n1708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1672  ( .A(\U1/aes_core/SB2/n1700 ), .B(
        \U1/aes_core/SB2/n1708 ), .Y(\U1/aes_core/SB2/n3248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1671  ( .A(\U1/aes_core/SB2/n3096 ), .B(
        \U1/aes_core/SB2/n3248 ), .Y(\U1/aes_core/SB2/n2987 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1670  ( .A(\U1/aes_core/SB2/n1203 ), .B(
        \U1/aes_core/SB2/n1158 ), .Y(\U1/aes_core/SB2/n1699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1669  ( .A(\U1/aes_core/SB2/n1690 ), .B(
        \U1/aes_core/SB2/n1699 ), .Y(\U1/aes_core/SB2/n3223 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1668  ( .A(\U1/aes_core/SB2/n3223 ), .Y(
        \U1/aes_core/SB2/n2968 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1667  ( .A0(\U1/aes_core/SB2/n3194 ), 
        .A1(\U1/aes_core/SB2/n2987 ), .B0(\U1/aes_core/SB2/n2968 ), .B1(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n1218 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1666  ( .AN(\U1/aes_core/SB2/n3009 ), 
        .B(\U1/aes_core/SB2/n1621 ), .C(\U1/aes_core/SB2/n1218 ), .Y(
        \U1/aes_core/SB2/n1721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1665  ( .A(\U1/aes_core/SB2/n1682 ), .B(
        \U1/aes_core/SB2/n1699 ), .Y(\U1/aes_core/SB2/n3113 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1664  ( .A(\U1/aes_core/SB2/n1686 ), .B(
        \U1/aes_core/SB2/n1687 ), .Y(\U1/aes_core/SB2/n3258 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1663  ( .A(\U1/aes_core/SB2/n1709 ), .B(
        \U1/aes_core/SB2/n1690 ), .Y(\U1/aes_core/SB2/n3164 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1662  ( .A(\U1/aes_core/SB2/n1686 ), .B(
        \U1/aes_core/SB2/n1692 ), .Y(\U1/aes_core/SB2/n3161 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1661  ( .A(\U1/aes_core/SB2/n1683 ), .B(
        \U1/aes_core/SB2/n1693 ), .Y(\U1/aes_core/SB2/n3166 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1660  ( .A(\U1/aes_core/SB2/n3166 ), .Y(
        \U1/aes_core/SB2/n3146 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1659  ( .A(\U1/aes_core/SB2/n3248 ), .Y(
        \U1/aes_core/SB2/n2982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1658  ( .A(\U1/aes_core/SB2/n1684 ), .B(
        \U1/aes_core/SB2/n1692 ), .Y(\U1/aes_core/SB2/n3184 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1657  ( .A(\U1/aes_core/SB2/n3184 ), .Y(
        \U1/aes_core/SB2/n3209 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1656  ( .A0(\U1/aes_core/SB2/n3146 ), 
        .A1(\U1/aes_core/SB2/n3210 ), .B0(\U1/aes_core/SB2/n2982 ), .B1(
        \U1/aes_core/SB2/n3209 ), .Y(\U1/aes_core/SB2/n1685 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1655  ( .A0(\U1/aes_core/SB2/n3113 ), 
        .A1(\U1/aes_core/SB2/n3258 ), .B0(\U1/aes_core/SB2/n3164 ), .B1(
        \U1/aes_core/SB2/n3161 ), .C0(\U1/aes_core/SB2/n1685 ), .Y(
        \U1/aes_core/SB2/n1720 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1654  ( .A(\U1/aes_core/SB2/n3166 ), .B(
        \U1/aes_core/SB2/n3113 ), .Y(\U1/aes_core/SB2/n2975 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1653  ( .A(\U1/aes_core/SB2/n3161 ), .B(
        \U1/aes_core/SB2/n3096 ), .Y(\U1/aes_core/SB2/n2985 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1652  ( .A(\U1/aes_core/SB2/n2985 ), .Y(
        \U1/aes_core/SB2/n1689 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1651  ( .A(\U1/aes_core/SB2/n1686 ), .B(
        \U1/aes_core/SB2/n1702 ), .Y(\U1/aes_core/SB2/n3236 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1650  ( .A(\U1/aes_core/SB2/n3236 ), .Y(
        \U1/aes_core/SB2/n3185 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1649  ( .A(\U1/aes_core/SB2/n1687 ), .B(
        \U1/aes_core/SB2/n1693 ), .Y(\U1/aes_core/SB2/n3221 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1648  ( .A(\U1/aes_core/SB2/n3221 ), .Y(
        \U1/aes_core/SB2/n3232 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1647  ( .A0(\U1/aes_core/SB2/n3185 ), 
        .A1(\U1/aes_core/SB2/n3232 ), .B0(\U1/aes_core/SB2/n3186 ), .Y(
        \U1/aes_core/SB2/n1688 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1646  ( .A(\U1/aes_core/SB2/n1691 ), .B(
        \U1/aes_core/SB2/n1708 ), .Y(\U1/aes_core/SB2/n3237 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1645  ( .A(\U1/aes_core/SB2/n3237 ), .Y(
        \U1/aes_core/SB2/n3187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1644  ( .A(\U1/aes_core/SB2/n3187 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3002 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1643  ( .AN(\U1/aes_core/SB2/n2975 ), 
        .B(\U1/aes_core/SB2/n1689 ), .C(\U1/aes_core/SB2/n1688 ), .D(
        \U1/aes_core/SB2/n3002 ), .Y(\U1/aes_core/SB2/n1698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1642  ( .A(\U1/aes_core/SB2/n1701 ), .B(
        \U1/aes_core/SB2/n1699 ), .Y(\U1/aes_core/SB2/n3257 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1641  ( .A(\U1/aes_core/SB2/n1691 ), .B(
        \U1/aes_core/SB2/n1690 ), .Y(\U1/aes_core/SB2/n3249 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1640  ( .A0(\U1/aes_core/SB2/n2327 ), 
        .A1(\U1/aes_core/SB2/n3076 ), .B0(\U1/aes_core/SB2/n3257 ), .B1(
        \U1/aes_core/SB2/n3166 ), .C0(\U1/aes_core/SB2/n3249 ), .C1(
        \U1/aes_core/SB2/n3184 ), .Y(\U1/aes_core/SB2/n1697 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1639  ( .A(\U1/aes_core/SB2/n3208 ), .B(
        \U1/aes_core/SB2/n2327 ), .Y(\U1/aes_core/SB2/n3060 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1638  ( .A(\U1/aes_core/SB2/n2982 ), .B(
        \U1/aes_core/SB2/n3146 ), .Y(\U1/aes_core/SB2/n3013 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1637  ( .A(\U1/aes_core/SB2/n3209 ), .B(
        \U1/aes_core/SB2/n3210 ), .Y(\U1/aes_core/SB2/n3033 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1636  ( .A(\U1/aes_core/SB2/n3164 ), .Y(
        \U1/aes_core/SB2/n3238 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1635  ( .A(\U1/aes_core/SB2/n3238 ), .B(
        \U1/aes_core/SB2/n3068 ), .Y(\U1/aes_core/SB2/n3071 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1634  ( .AN(\U1/aes_core/SB2/n3060 ), 
        .B(\U1/aes_core/SB2/n3013 ), .C(\U1/aes_core/SB2/n3033 ), .D(
        \U1/aes_core/SB2/n3071 ), .Y(\U1/aes_core/SB2/n1696 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1633  ( .A(\U1/aes_core/SB2/n1709 ), .B(
        \U1/aes_core/SB2/n1701 ), .Y(\U1/aes_core/SB2/n2983 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1632  ( .A(\U1/aes_core/SB2/n2983 ), .B(
        \U1/aes_core/SB2/n3220 ), .Y(\U1/aes_core/SB2/n3137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1631  ( .A(\U1/aes_core/SB2/n1693 ), .B(
        \U1/aes_core/SB2/n1692 ), .Y(\U1/aes_core/SB2/n3256 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1630  ( .A(\U1/aes_core/SB2/n3223 ), .B(
        \U1/aes_core/SB2/n3256 ), .Y(\U1/aes_core/SB2/n3102 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1629  ( .A(\U1/aes_core/SB2/n3102 ), .Y(
        \U1/aes_core/SB2/n1694 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1628  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3068 ), .Y(\U1/aes_core/SB2/n3121 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1627  ( .A(\U1/aes_core/SB2/n3256 ), .Y(
        \U1/aes_core/SB2/n3239 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1626  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3239 ), .Y(\U1/aes_core/SB2/n3172 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1625  ( .AN(\U1/aes_core/SB2/n3137 ), 
        .B(\U1/aes_core/SB2/n1694 ), .C(\U1/aes_core/SB2/n3121 ), .D(
        \U1/aes_core/SB2/n3172 ), .Y(\U1/aes_core/SB2/n1695 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1624  ( .A(\U1/aes_core/SB2/n1698 ), .B(
        \U1/aes_core/SB2/n1697 ), .C(\U1/aes_core/SB2/n1696 ), .D(
        \U1/aes_core/SB2/n1695 ), .Y(\U1/aes_core/SB2/n2905 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1623  ( .A(\U1/aes_core/SB2/n3163 ), .B(
        \U1/aes_core/SB2/n2983 ), .Y(\U1/aes_core/SB2/n3171 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1622  ( .A(\U1/aes_core/SB2/n1708 ), .B(
        \U1/aes_core/SB2/n1699 ), .Y(\U1/aes_core/SB2/n3079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1621  ( .A(\U1/aes_core/SB2/n3145 ), .B(
        \U1/aes_core/SB2/n3079 ), .Y(\U1/aes_core/SB2/n3050 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1620  ( .A(\U1/aes_core/SB2/n3257 ), .Y(
        \U1/aes_core/SB2/n3213 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1619  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3194 ), .Y(\U1/aes_core/SB2/n2999 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1618  ( .A0(\U1/aes_core/SB2/n3079 ), 
        .A1(\U1/aes_core/SB2/n3256 ), .B0(\U1/aes_core/SB2/n2999 ), .Y(
        \U1/aes_core/SB2/n1707 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1617  ( .A(\U1/aes_core/SB2/n3094 ), .Y(
        \U1/aes_core/SB2/n3189 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1616  ( .A(\U1/aes_core/SB2/n3189 ), .B(
        \U1/aes_core/SB2/n3212 ), .Y(\U1/aes_core/SB2/n3190 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1615  ( .A(\U1/aes_core/SB2/n3212 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1614  ( .A(\U1/aes_core/SB2/n1701 ), .B(
        \U1/aes_core/SB2/n1700 ), .Y(\U1/aes_core/SB2/n3219 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1613  ( .A(\U1/aes_core/SB2/n3219 ), .Y(
        \U1/aes_core/SB2/n2994 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1612  ( .A(\U1/aes_core/SB2/n3185 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3018 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1611  ( .A(\U1/aes_core/SB2/n3207 ), .Y(
        \U1/aes_core/SB2/n3188 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1610  ( .A(\U1/aes_core/SB2/n3188 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3082 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1609  ( .A(\U1/aes_core/SB2/n3190 ), .B(
        \U1/aes_core/SB2/n3149 ), .C(\U1/aes_core/SB2/n3018 ), .D(
        \U1/aes_core/SB2/n3082 ), .Y(\U1/aes_core/SB2/n1706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1608  ( .A(\U1/aes_core/SB2/n3209 ), .B(
        \U1/aes_core/SB2/n3187 ), .Y(\U1/aes_core/SB2/n3116 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1607  ( .A(\U1/aes_core/SB2/n3251 ), .B(
        \U1/aes_core/SB2/n3187 ), .Y(\U1/aes_core/SB2/n3107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1606  ( .A(\U1/aes_core/SB2/n3249 ), .Y(
        \U1/aes_core/SB2/n3242 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1605  ( .A(\U1/aes_core/SB2/n3146 ), .B(
        \U1/aes_core/SB2/n3242 ), .Y(\U1/aes_core/SB2/n2979 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1604  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3185 ), .Y(\U1/aes_core/SB2/n3090 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1603  ( .A(\U1/aes_core/SB2/n3116 ), .B(
        \U1/aes_core/SB2/n3107 ), .C(\U1/aes_core/SB2/n2979 ), .D(
        \U1/aes_core/SB2/n3090 ), .Y(\U1/aes_core/SB2/n1705 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1602  ( .A(\U1/aes_core/SB2/n3161 ), .Y(
        \U1/aes_core/SB2/n3130 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1601  ( .A(\U1/aes_core/SB2/n2982 ), .B(
        \U1/aes_core/SB2/n3130 ), .Y(\U1/aes_core/SB2/n2966 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1600  ( .A(\U1/aes_core/SB2/n1703 ), .B(
        \U1/aes_core/SB2/n1702 ), .Y(\U1/aes_core/SB2/n3196 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1599  ( .A(\U1/aes_core/SB2/n3196 ), .Y(
        \U1/aes_core/SB2/n3230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1598  ( .A(\U1/aes_core/SB2/n2982 ), .B(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n3030 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1597  ( .A(\U1/aes_core/SB2/n3145 ), .Y(
        \U1/aes_core/SB2/n3253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1596  ( .A(\U1/aes_core/SB2/n3253 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n3065 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1595  ( .A(\U1/aes_core/SB2/n3186 ), .B(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n3214 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1594  ( .A(\U1/aes_core/SB2/n2966 ), .B(
        \U1/aes_core/SB2/n3030 ), .C(\U1/aes_core/SB2/n3065 ), .D(
        \U1/aes_core/SB2/n3214 ), .Y(\U1/aes_core/SB2/n1704 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1593  ( .A(\U1/aes_core/SB2/n3171 ), .B(
        \U1/aes_core/SB2/n3050 ), .C(\U1/aes_core/SB2/n1707 ), .D(
        \U1/aes_core/SB2/n1706 ), .E(\U1/aes_core/SB2/n1705 ), .F(
        \U1/aes_core/SB2/n1704 ), .Y(\U1/aes_core/SB2/n2894 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1592  ( .A(\U1/aes_core/SB2/n2894 ), .Y(
        \U1/aes_core/SB2/n1718 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1591  ( .A(\U1/aes_core/SB2/n3221 ), .B(
        \U1/aes_core/SB2/n3079 ), .Y(\U1/aes_core/SB2/n2976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1590  ( .A(\U1/aes_core/SB2/n1709 ), .B(
        \U1/aes_core/SB2/n1708 ), .Y(\U1/aes_core/SB2/n3218 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1589  ( .A(\U1/aes_core/SB2/n3218 ), .B(
        \U1/aes_core/SB2/n3094 ), .Y(\U1/aes_core/SB2/n3103 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1588  ( .A(\U1/aes_core/SB2/n3103 ), .Y(
        \U1/aes_core/SB2/n1711 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1587  ( .A(\U1/aes_core/SB2/n3096 ), .Y(
        \U1/aes_core/SB2/n3243 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1586  ( .A0(\U1/aes_core/SB2/n2994 ), 
        .A1(\U1/aes_core/SB2/n3243 ), .B0(\U1/aes_core/SB2/n3230 ), .Y(
        \U1/aes_core/SB2/n1710 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1585  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3130 ), .Y(\U1/aes_core/SB2/n3001 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1584  ( .AN(\U1/aes_core/SB2/n2976 ), 
        .B(\U1/aes_core/SB2/n1711 ), .C(\U1/aes_core/SB2/n1710 ), .D(
        \U1/aes_core/SB2/n3001 ), .Y(\U1/aes_core/SB2/n1715 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1583  ( .A0(\U1/aes_core/SB2/n3207 ), 
        .A1(\U1/aes_core/SB2/n3255 ), .B0(\U1/aes_core/SB2/n3113 ), .B1(
        \U1/aes_core/SB2/n3161 ), .C0(\U1/aes_core/SB2/n3220 ), .C1(
        \U1/aes_core/SB2/n3237 ), .Y(\U1/aes_core/SB2/n1714 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1582  ( .A(\U1/aes_core/SB2/n3255 ), .B(
        \U1/aes_core/SB2/n3258 ), .Y(\U1/aes_core/SB2/n3041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1581  ( .A(\U1/aes_core/SB2/n3243 ), .B(
        \U1/aes_core/SB2/n3185 ), .Y(\U1/aes_core/SB2/n3174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1580  ( .A(\U1/aes_core/SB2/n3146 ), .B(
        \U1/aes_core/SB2/n3243 ), .Y(\U1/aes_core/SB2/n3108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1579  ( .A(\U1/aes_core/SB2/n3130 ), .B(
        \U1/aes_core/SB2/n3210 ), .Y(\U1/aes_core/SB2/n2980 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1578  ( .AN(\U1/aes_core/SB2/n3041 ), 
        .B(\U1/aes_core/SB2/n3174 ), .C(\U1/aes_core/SB2/n3108 ), .D(
        \U1/aes_core/SB2/n2980 ), .Y(\U1/aes_core/SB2/n1713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1577  ( .A(\U1/aes_core/SB2/n3253 ), .B(
        \U1/aes_core/SB2/n3238 ), .Y(\U1/aes_core/SB2/n3053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1576  ( .A(\U1/aes_core/SB2/n3130 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3120 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1575  ( .A(\U1/aes_core/SB2/n2982 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3021 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1574  ( .A(\U1/aes_core/SB2/n3189 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n3066 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1573  ( .A(\U1/aes_core/SB2/n3053 ), .B(
        \U1/aes_core/SB2/n3120 ), .C(\U1/aes_core/SB2/n3021 ), .D(
        \U1/aes_core/SB2/n3066 ), .Y(\U1/aes_core/SB2/n1712 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1572  ( .A(\U1/aes_core/SB2/n1715 ), .B(
        \U1/aes_core/SB2/n1714 ), .C(\U1/aes_core/SB2/n1713 ), .D(
        \U1/aes_core/SB2/n1712 ), .Y(\U1/aes_core/SB2/n1716 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1571  ( .A(\U1/aes_core/SB2/n1716 ), .Y(
        \U1/aes_core/SB2/n3235 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1570  ( .A(\U1/aes_core/SB2/n3251 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n1717 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1569  ( .AN(\U1/aes_core/SB2/n2905 ), 
        .B(\U1/aes_core/SB2/n1718 ), .C(\U1/aes_core/SB2/n3235 ), .D(
        \U1/aes_core/SB2/n1717 ), .Y(\U1/aes_core/SB2/n1719 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1568  ( .A(\U1/aes_core/SB2/n3014 ), .B(
        \U1/aes_core/SB2/n3111 ), .C(\U1/aes_core/SB2/n1722 ), .D(
        \U1/aes_core/SB2/n1721 ), .E(\U1/aes_core/SB2/n1720 ), .F(
        \U1/aes_core/SB2/n1719 ), .Y(\U1/aes_core/SB2/n2346 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1567  ( .A(\U1/aes_core/SB2/n3236 ), .B(
        \U1/aes_core/SB2/n2327 ), .Y(\U1/aes_core/SB2/n3059 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1566  ( .A(\U1/aes_core/SB2/n3186 ), .B(
        \U1/aes_core/SB2/n3253 ), .Y(\U1/aes_core/SB2/n3110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1565  ( .A(\U1/aes_core/SB2/n3242 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3012 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1564  ( .A(\U1/aes_core/SB2/n2983 ), .Y(
        \U1/aes_core/SB2/n3231 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1563  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3035 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1562  ( .AN(\U1/aes_core/SB2/n3059 ), 
        .B(\U1/aes_core/SB2/n3110 ), .C(\U1/aes_core/SB2/n3012 ), .D(
        \U1/aes_core/SB2/n3035 ), .Y(\U1/aes_core/SB2/n1729 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1561  ( .A(\U1/aes_core/SB2/n3223 ), .B(
        \U1/aes_core/SB2/n3094 ), .Y(\U1/aes_core/SB2/n3136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1560  ( .A(\U1/aes_core/SB2/n3146 ), .B(
        \U1/aes_core/SB2/n3212 ), .Y(\U1/aes_core/SB2/n2992 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1559  ( .A0(\U1/aes_core/SB2/n3232 ), 
        .A1(\U1/aes_core/SB2/n3152 ), .B0(\U1/aes_core/SB2/n2982 ), .Y(
        \U1/aes_core/SB2/n1723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1558  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3084 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1557  ( .AN(\U1/aes_core/SB2/n3136 ), 
        .B(\U1/aes_core/SB2/n2992 ), .C(\U1/aes_core/SB2/n1723 ), .D(
        \U1/aes_core/SB2/n3084 ), .Y(\U1/aes_core/SB2/n1724 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1556  ( .A(\U1/aes_core/SB2/n1724 ), .Y(
        \U1/aes_core/SB2/n1728 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1555  ( .A(\U1/aes_core/SB2/n3113 ), .Y(
        \U1/aes_core/SB2/n3233 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1554  ( .A(\U1/aes_core/SB2/n3258 ), .Y(
        \U1/aes_core/SB2/n3153 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U1553  ( .A0(\U1/aes_core/SB2/n3253 ), 
        .A1(\U1/aes_core/SB2/n3187 ), .B0(\U1/aes_core/SB2/n3233 ), .B1(
        \U1/aes_core/SB2/n3068 ), .C0(\U1/aes_core/SB2/n3153 ), .C1(
        \U1/aes_core/SB2/n3231 ), .Y(\U1/aes_core/SB2/n1727 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1552  ( .A0(\U1/aes_core/SB2/n3079 ), 
        .A1(\U1/aes_core/SB2/n3236 ), .B0(\U1/aes_core/SB2/n3256 ), .B1(
        \U1/aes_core/SB2/n3257 ), .Y(\U1/aes_core/SB2/n1725 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1551  ( .A0(\U1/aes_core/SB2/n3130 ), 
        .A1(\U1/aes_core/SB2/n2968 ), .B0(\U1/aes_core/SB2/n3186 ), .B1(
        \U1/aes_core/SB2/n3209 ), .C0(\U1/aes_core/SB2/n1725 ), .Y(
        \U1/aes_core/SB2/n1726 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1550  ( .AN(\U1/aes_core/SB2/n1729 ), 
        .B(\U1/aes_core/SB2/n1728 ), .C(\U1/aes_core/SB2/n1727 ), .D(
        \U1/aes_core/SB2/n1726 ), .Y(\U1/aes_core/SB2/n2903 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1549  ( .A(\U1/aes_core/SB2/n3257 ), .B(
        \U1/aes_core/SB2/n3094 ), .Y(\U1/aes_core/SB2/n2977 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1548  ( .A0(\U1/aes_core/SB2/n3164 ), 
        .A1(\U1/aes_core/SB2/n3257 ), .B0(\U1/aes_core/SB2/n3196 ), .Y(
        \U1/aes_core/SB2/n1734 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1547  ( .A(\U1/aes_core/SB2/n3196 ), .B(
        \U1/aes_core/SB2/n3184 ), .Y(\U1/aes_core/SB2/n3061 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB2/U1546  ( .A0(\U1/aes_core/SB2/n3185 ), 
        .A1(\U1/aes_core/SB2/n2968 ), .B0(\U1/aes_core/SB2/n3061 ), .B1(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n1733 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1545  ( .A0(\U1/aes_core/SB2/n3218 ), 
        .A1(\U1/aes_core/SB2/n3258 ), .B0(\U1/aes_core/SB2/n2983 ), .B1(
        \U1/aes_core/SB2/n3076 ), .C0(\U1/aes_core/SB2/n3220 ), .C1(
        \U1/aes_core/SB2/n3249 ), .Y(\U1/aes_core/SB2/n1732 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1544  ( .A(\U1/aes_core/SB2/n3079 ), .Y(
        \U1/aes_core/SB2/n3147 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1543  ( .A(\U1/aes_core/SB2/n3251 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3173 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1542  ( .A(\U1/aes_core/SB2/n3146 ), .B(
        \U1/aes_core/SB2/n2968 ), .Y(\U1/aes_core/SB2/n3000 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1541  ( .A(\U1/aes_core/SB2/n2982 ), .B(
        \U1/aes_core/SB2/n3189 ), .Y(\U1/aes_core/SB2/n3020 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1540  ( .A(\U1/aes_core/SB2/n3146 ), .B(
        \U1/aes_core/SB2/n3187 ), .Y(\U1/aes_core/SB2/n3119 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1539  ( .A(\U1/aes_core/SB2/n3173 ), .B(
        \U1/aes_core/SB2/n3000 ), .C(\U1/aes_core/SB2/n3020 ), .D(
        \U1/aes_core/SB2/n3119 ), .Y(\U1/aes_core/SB2/n1731 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1538  ( .A(\U1/aes_core/SB2/n3166 ), .B(
        \U1/aes_core/SB2/n3079 ), .Y(\U1/aes_core/SB2/n3042 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1537  ( .A(\U1/aes_core/SB2/n3152 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3052 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1536  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3068 ), .Y(\U1/aes_core/SB2/n3083 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1535  ( .AN(\U1/aes_core/SB2/n3042 ), 
        .B(\U1/aes_core/SB2/n3052 ), .C(\U1/aes_core/SB2/n3083 ), .Y(
        \U1/aes_core/SB2/n1730 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1534  ( .A(\U1/aes_core/SB2/n2977 ), .B(
        \U1/aes_core/SB2/n1734 ), .C(\U1/aes_core/SB2/n1733 ), .D(
        \U1/aes_core/SB2/n1732 ), .E(\U1/aes_core/SB2/n1731 ), .F(
        \U1/aes_core/SB2/n1730 ), .Y(\U1/aes_core/SB2/n3264 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1533  ( .A0(\U1/aes_core/SB2/n2982 ), 
        .A1(\U1/aes_core/SB2/n3210 ), .B0(\U1/aes_core/SB2/n3241 ), .Y(
        \U1/aes_core/SB2/n1735 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1532  ( .A(\U1/aes_core/SB2/n2968 ), .B(
        \U1/aes_core/SB2/n3068 ), .Y(\U1/aes_core/SB2/n3105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1531  ( .A(\U1/aes_core/SB2/n3185 ), .B(
        \U1/aes_core/SB2/n3233 ), .Y(\U1/aes_core/SB2/n2997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1530  ( .A(\U1/aes_core/SB2/n3233 ), .B(
        \U1/aes_core/SB2/n3189 ), .Y(\U1/aes_core/SB2/n3048 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1529  ( .A(\U1/aes_core/SB2/n1735 ), .B(
        \U1/aes_core/SB2/n3105 ), .C(\U1/aes_core/SB2/n2997 ), .D(
        \U1/aes_core/SB2/n3048 ), .Y(\U1/aes_core/SB2/n1739 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1528  ( .A0(\U1/aes_core/SB2/n3236 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n2983 ), .B1(
        \U1/aes_core/SB2/n3208 ), .C0(\U1/aes_core/SB2/n3237 ), .C1(
        \U1/aes_core/SB2/n3094 ), .Y(\U1/aes_core/SB2/n1738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1527  ( .A(\U1/aes_core/SB2/n3188 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n3029 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1526  ( .A(\U1/aes_core/SB2/n3187 ), .B(
        \U1/aes_core/SB2/n3239 ), .Y(\U1/aes_core/SB2/n3169 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1525  ( .A(\U1/aes_core/SB2/n3187 ), .B(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n3016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1524  ( .A(\U1/aes_core/SB2/n3242 ), .B(
        \U1/aes_core/SB2/n3232 ), .Y(\U1/aes_core/SB2/n2978 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1523  ( .A(\U1/aes_core/SB2/n3029 ), .B(
        \U1/aes_core/SB2/n3169 ), .C(\U1/aes_core/SB2/n3016 ), .D(
        \U1/aes_core/SB2/n2978 ), .Y(\U1/aes_core/SB2/n1737 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1522  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1521  ( .A(\U1/aes_core/SB2/n3251 ), .B(
        \U1/aes_core/SB2/n3212 ), .Y(\U1/aes_core/SB2/n3064 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1520  ( .A(\U1/aes_core/SB2/n3241 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1519  ( .A(\U1/aes_core/SB2/n2994 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n2965 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1518  ( .A(\U1/aes_core/SB2/n3091 ), .B(
        \U1/aes_core/SB2/n3064 ), .C(\U1/aes_core/SB2/n3115 ), .D(
        \U1/aes_core/SB2/n2965 ), .Y(\U1/aes_core/SB2/n1736 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1517  ( .A(\U1/aes_core/SB2/n1739 ), .B(
        \U1/aes_core/SB2/n1738 ), .C(\U1/aes_core/SB2/n1737 ), .D(
        \U1/aes_core/SB2/n1736 ), .Y(\U1/aes_core/SB2/n2892 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1516  ( .A(\U1/aes_core/SB2/n2346 ), .B(
        \U1/aes_core/SB2/n2903 ), .C(\U1/aes_core/SB2/n3264 ), .D(
        \U1/aes_core/SB2/n2892 ), .Y(\U1/aes_core/SB2/n1748 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1515  ( .A(\U1/aes_core/SB2/n3218 ), .Y(
        \U1/aes_core/SB2/n3142 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1514  ( .A0(\U1/aes_core/SB2/n3094 ), 
        .A1(\U1/aes_core/SB2/n2328 ), .B0(\U1/aes_core/SB2/n3063 ), .B1(
        \U1/aes_core/SB2/n3249 ), .Y(\U1/aes_core/SB2/n1740 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1513  ( .A0(\U1/aes_core/SB2/n3142 ), 
        .A1(\U1/aes_core/SB2/n3194 ), .B0(\U1/aes_core/SB2/n3243 ), .B1(
        \U1/aes_core/SB2/n3251 ), .C0(\U1/aes_core/SB2/n1740 ), .Y(
        \U1/aes_core/SB2/n1747 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1512  ( .A(\U1/aes_core/SB2/n3163 ), .B(
        \U1/aes_core/SB2/n3166 ), .Y(\U1/aes_core/SB2/n3162 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1511  ( .A0(\U1/aes_core/SB2/n3097 ), 
        .A1(\U1/aes_core/SB2/n3166 ), .B0(\U1/aes_core/SB2/n3079 ), .B1(
        \U1/aes_core/SB2/n3207 ), .Y(\U1/aes_core/SB2/n1741 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1510  ( .A0(\U1/aes_core/SB2/n2994 ), 
        .A1(\U1/aes_core/SB2/n3162 ), .B0(\U1/aes_core/SB2/n3213 ), .B1(
        \U1/aes_core/SB2/n3232 ), .C0(\U1/aes_core/SB2/n1741 ), .Y(
        \U1/aes_core/SB2/n1746 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1509  ( .A(\U1/aes_core/SB2/n3237 ), .B(
        \U1/aes_core/SB2/n3096 ), .Y(\U1/aes_core/SB2/n1744 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1508  ( .A(\U1/aes_core/SB2/n3187 ), .B(
        \U1/aes_core/SB2/n3212 ), .Y(\U1/aes_core/SB2/n3154 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1507  ( .A(\U1/aes_core/SB2/n3154 ), .Y(
        \U1/aes_core/SB2/n1743 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1506  ( .A(\U1/aes_core/SB2/n3145 ), .B(
        \U1/aes_core/SB2/n3218 ), .Y(\U1/aes_core/SB2/n3026 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1505  ( .A(\U1/aes_core/SB2/n3223 ), .B(
        \U1/aes_core/SB2/n3221 ), .Y(\U1/aes_core/SB2/n3179 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1503  ( .A(\U1/aes_core/SB2/n3194 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3036 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1501  ( .A0(\U1/aes_core/SB2/n3153 ), 
        .A1(\U1/aes_core/SB2/n1744 ), .B0(\U1/aes_core/SB2/n3130 ), .B1(
        \U1/aes_core/SB2/n1743 ), .C0(\U1/aes_core/SB2/n1742 ), .Y(
        \U1/aes_core/SB2/n1745 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1500  ( .AN(\U1/aes_core/SB2/n1748 ), 
        .B(\U1/aes_core/SB2/n1747 ), .C(\U1/aes_core/SB2/n1746 ), .D(
        \U1/aes_core/SB2/n1745 ), .Y(\U1/aes_core/sb2 [0]) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1499  ( .A(Dout[46]), .Y(
        \U1/aes_core/SB2/n1755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1498  ( .A(Dout[47]), .Y(
        \U1/aes_core/SB2/n1750 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1497  ( .A(\U1/aes_core/SB2/n1755 ), .B(
        \U1/aes_core/SB2/n1750 ), .Y(\U1/aes_core/SB2/n1760 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1496  ( .A(Dout[45]), .Y(
        \U1/aes_core/SB2/n1749 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1495  ( .A(\U1/aes_core/SB2/n1749 ), .B(
        Dout[44]), .Y(\U1/aes_core/SB2/n1767 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1494  ( .A(\U1/aes_core/SB2/n1760 ), .B(
        \U1/aes_core/SB2/n1767 ), .Y(\U1/aes_core/SB2/n3300 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1493  ( .A(Dout[43]), .Y(
        \U1/aes_core/SB2/n1758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1492  ( .A(\U1/aes_core/SB2/n1758 ), .B(
        Dout[42]), .Y(\U1/aes_core/SB2/n1773 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1491  ( .A(Dout[40]), .Y(
        \U1/aes_core/SB2/n1751 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1490  ( .A(\U1/aes_core/SB2/n1751 ), .B(
        Dout[41]), .Y(\U1/aes_core/SB2/n1761 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1489  ( .A(\U1/aes_core/SB2/n1773 ), .B(
        \U1/aes_core/SB2/n1761 ), .Y(\U1/aes_core/SB2/n1912 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1488  ( .A(\U1/aes_core/SB2/n3300 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n1821 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1487  ( .A(Dout[41]), .Y(
        \U1/aes_core/SB2/n1752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1486  ( .A(\U1/aes_core/SB2/n1752 ), .B(
        Dout[40]), .Y(\U1/aes_core/SB2/n1770 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1485  ( .A(Dout[42]), .Y(
        \U1/aes_core/SB2/n1757 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1484  ( .A(\U1/aes_core/SB2/n1757 ), .B(
        Dout[43]), .Y(\U1/aes_core/SB2/n1754 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1483  ( .A(\U1/aes_core/SB2/n1770 ), .B(
        \U1/aes_core/SB2/n1754 ), .Y(\U1/aes_core/SB2/n3346 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1482  ( .A(Dout[44]), .Y(
        \U1/aes_core/SB2/n1753 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1481  ( .A(\U1/aes_core/SB2/n1749 ), .B(
        \U1/aes_core/SB2/n1753 ), .Y(\U1/aes_core/SB2/n1781 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1480  ( .A(\U1/aes_core/SB2/n1750 ), .B(
        Dout[46]), .Y(\U1/aes_core/SB2/n1756 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1479  ( .A(\U1/aes_core/SB2/n1781 ), .B(
        \U1/aes_core/SB2/n1756 ), .Y(\U1/aes_core/SB2/n2021 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1478  ( .A0(\U1/aes_core/SB2/n1912 ), 
        .A1(\U1/aes_core/SB2/n3346 ), .B0(\U1/aes_core/SB2/n2021 ), .Y(
        \U1/aes_core/SB2/n1766 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1477  ( .A(\U1/aes_core/SB2/n1752 ), .B(
        \U1/aes_core/SB2/n1751 ), .Y(\U1/aes_core/SB2/n1772 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1476  ( .A(\U1/aes_core/SB2/n1754 ), .B(
        \U1/aes_core/SB2/n1772 ), .Y(\U1/aes_core/SB2/n2020 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1475  ( .A(\U1/aes_core/SB2/n1753 ), .B(
        Dout[45]), .Y(\U1/aes_core/SB2/n1783 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1474  ( .A(\U1/aes_core/SB2/n1760 ), .B(
        \U1/aes_core/SB2/n1783 ), .Y(\U1/aes_core/SB2/n1995 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1473  ( .A(Dout[43]), .B(Dout[42]), .Y(
        \U1/aes_core/SB2/n1780 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1472  ( .A(\U1/aes_core/SB2/n1772 ), .B(
        \U1/aes_core/SB2/n1780 ), .Y(\U1/aes_core/SB2/n3301 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1471  ( .A(\U1/aes_core/SB2/n3301 ), .Y(
        \U1/aes_core/SB2/n3339 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1470  ( .A(Dout[41]), .B(Dout[40]), .Y(
        \U1/aes_core/SB2/n1779 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1469  ( .A(\U1/aes_core/SB2/n1754 ), .B(
        \U1/aes_core/SB2/n1779 ), .Y(\U1/aes_core/SB2/n3296 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1468  ( .A(\U1/aes_core/SB2/n3296 ), .Y(
        \U1/aes_core/SB2/n3333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1467  ( .A(\U1/aes_core/SB2/n3339 ), .B(
        \U1/aes_core/SB2/n3333 ), .Y(\U1/aes_core/SB2/n1823 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1466  ( .A(Dout[47]), .B(Dout[46]), .Y(
        \U1/aes_core/SB2/n1774 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1465  ( .A(\U1/aes_core/SB2/n1767 ), .B(
        \U1/aes_core/SB2/n1774 ), .Y(\U1/aes_core/SB2/n3309 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1464  ( .A0(\U1/aes_core/SB2/n2020 ), 
        .A1(\U1/aes_core/SB2/n1995 ), .B0(\U1/aes_core/SB2/n1823 ), .B1(
        \U1/aes_core/SB2/n3309 ), .Y(\U1/aes_core/SB2/n1765 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1463  ( .A(\U1/aes_core/SB2/n1754 ), .B(
        \U1/aes_core/SB2/n1761 ), .Y(\U1/aes_core/SB2/n1888 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1462  ( .A(\U1/aes_core/SB2/n1767 ), .B(
        \U1/aes_core/SB2/n1756 ), .Y(\U1/aes_core/SB2/n3344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1461  ( .A(Dout[45]), .B(Dout[44]), .Y(
        \U1/aes_core/SB2/n1759 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1460  ( .A(\U1/aes_core/SB2/n1760 ), .B(
        \U1/aes_core/SB2/n1759 ), .Y(\U1/aes_core/SB2/n3280 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1459  ( .A(\U1/aes_core/SB2/n1783 ), .B(
        \U1/aes_core/SB2/n1756 ), .Y(\U1/aes_core/SB2/n3278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1458  ( .A(\U1/aes_core/SB2/n1773 ), .B(
        \U1/aes_core/SB2/n1779 ), .Y(\U1/aes_core/SB2/n2010 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1457  ( .A0(\U1/aes_core/SB2/n1888 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n3301 ), .B1(
        \U1/aes_core/SB2/n3280 ), .C0(\U1/aes_core/SB2/n3278 ), .C1(
        \U1/aes_core/SB2/n2010 ), .Y(\U1/aes_core/SB2/n1764 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1456  ( .A(\U1/aes_core/SB2/n1755 ), .B(
        Dout[47]), .Y(\U1/aes_core/SB2/n1782 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1455  ( .A(\U1/aes_core/SB2/n1782 ), .B(
        \U1/aes_core/SB2/n1759 ), .Y(\U1/aes_core/SB2/n3308 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1454  ( .A(\U1/aes_core/SB2/n3308 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n1873 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1453  ( .A(\U1/aes_core/SB2/n1770 ), .B(
        \U1/aes_core/SB2/n1773 ), .Y(\U1/aes_core/SB2/n3342 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1452  ( .A(\U1/aes_core/SB2/n3342 ), .Y(
        \U1/aes_core/SB2/n2058 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1451  ( .A(\U1/aes_core/SB2/n1759 ), .B(
        \U1/aes_core/SB2/n1756 ), .Y(\U1/aes_core/SB2/n1806 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1450  ( .A(\U1/aes_core/SB2/n1806 ), .Y(
        \U1/aes_core/SB2/n3268 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1449  ( .A(\U1/aes_core/SB2/n2058 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n1856 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1448  ( .A(\U1/aes_core/SB2/n1758 ), .B(
        \U1/aes_core/SB2/n1757 ), .Y(\U1/aes_core/SB2/n1769 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1447  ( .A(\U1/aes_core/SB2/n1772 ), .B(
        \U1/aes_core/SB2/n1769 ), .Y(\U1/aes_core/SB2/n2006 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1446  ( .A(\U1/aes_core/SB2/n2006 ), .Y(
        \U1/aes_core/SB2/n2068 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U1445  ( .A(\U1/aes_core/SB2/n1774 ), .B(
        \U1/aes_core/SB2/n1759 ), .Y(\U1/aes_core/SB2/n3299 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1444  ( .A(\U1/aes_core/SB2/n2068 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1928 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1443  ( .A(\U1/aes_core/SB2/n1760 ), .B(
        \U1/aes_core/SB2/n1781 ), .Y(\U1/aes_core/SB2/n3347 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1442  ( .A(\U1/aes_core/SB2/n3347 ), .Y(
        \U1/aes_core/SB2/n3305 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1441  ( .A(\U1/aes_core/SB2/n3305 ), .B(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n1953 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1440  ( .AN(\U1/aes_core/SB2/n1873 ), 
        .B(\U1/aes_core/SB2/n1856 ), .C(\U1/aes_core/SB2/n1928 ), .D(
        \U1/aes_core/SB2/n1953 ), .Y(\U1/aes_core/SB2/n1763 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1439  ( .A(\U1/aes_core/SB2/n1995 ), .Y(
        \U1/aes_core/SB2/n3269 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1438  ( .A(\U1/aes_core/SB2/n1780 ), .B(
        \U1/aes_core/SB2/n1761 ), .Y(\U1/aes_core/SB2/n2017 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1437  ( .A(\U1/aes_core/SB2/n2017 ), .Y(
        \U1/aes_core/SB2/n2054 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1436  ( .A(\U1/aes_core/SB2/n3269 ), .B(
        \U1/aes_core/SB2/n2054 ), .Y(\U1/aes_core/SB2/n1843 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1435  ( .A(\U1/aes_core/SB2/n3278 ), .Y(
        \U1/aes_core/SB2/n3332 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1434  ( .A(\U1/aes_core/SB2/n1761 ), .B(
        \U1/aes_core/SB2/n1769 ), .Y(\U1/aes_core/SB2/n2057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1433  ( .A(\U1/aes_core/SB2/n2057 ), .Y(
        \U1/aes_core/SB2/n2019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1432  ( .A(\U1/aes_core/SB2/n3332 ), .B(
        \U1/aes_core/SB2/n2019 ), .Y(\U1/aes_core/SB2/n1879 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1431  ( .A(\U1/aes_core/SB2/n3269 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1966 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U1430  ( .A(\U1/aes_core/SB2/n1843 ), .B(
        \U1/aes_core/SB2/n1879 ), .C(\U1/aes_core/SB2/n1966 ), .Y(
        \U1/aes_core/SB2/n1762 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1429  ( .A(\U1/aes_core/SB2/n1821 ), .B(
        \U1/aes_core/SB2/n1766 ), .C(\U1/aes_core/SB2/n1765 ), .D(
        \U1/aes_core/SB2/n1764 ), .E(\U1/aes_core/SB2/n1763 ), .F(
        \U1/aes_core/SB2/n1762 ), .Y(\U1/aes_core/SB2/n3353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1428  ( .A(\U1/aes_core/SB2/n1995 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n1944 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1427  ( .A(\U1/aes_core/SB2/n2010 ), .Y(
        \U1/aes_core/SB2/n3330 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1426  ( .A(\U1/aes_core/SB2/n1888 ), .Y(
        \U1/aes_core/SB2/n3334 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1425  ( .A(\U1/aes_core/SB2/n1767 ), .B(
        \U1/aes_core/SB2/n1782 ), .Y(\U1/aes_core/SB2/n3343 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1424  ( .A(\U1/aes_core/SB2/n3343 ), .Y(
        \U1/aes_core/SB2/n3274 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1423  ( .A0(\U1/aes_core/SB2/n3330 ), 
        .A1(\U1/aes_core/SB2/n3334 ), .B0(\U1/aes_core/SB2/n3274 ), .Y(
        \U1/aes_core/SB2/n1768 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1422  ( .A(\U1/aes_core/SB2/n3305 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1903 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1421  ( .A(\U1/aes_core/SB2/n2021 ), .Y(
        \U1/aes_core/SB2/n2053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1420  ( .A(\U1/aes_core/SB2/n3339 ), .B(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n1865 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1419  ( .AN(\U1/aes_core/SB2/n1944 ), 
        .B(\U1/aes_core/SB2/n1768 ), .C(\U1/aes_core/SB2/n1903 ), .D(
        \U1/aes_core/SB2/n1865 ), .Y(\U1/aes_core/SB2/n1778 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1418  ( .A(\U1/aes_core/SB2/n3309 ), .Y(
        \U1/aes_core/SB2/n1976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1417  ( .A(\U1/aes_core/SB2/n1770 ), .B(
        \U1/aes_core/SB2/n1780 ), .Y(\U1/aes_core/SB2/n2039 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1416  ( .A(\U1/aes_core/SB2/n2039 ), .Y(
        \U1/aes_core/SB2/n3340 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1415  ( .A(\U1/aes_core/SB2/n3280 ), .Y(
        \U1/aes_core/SB2/n2055 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1414  ( .A(\U1/aes_core/SB2/n1779 ), .B(
        \U1/aes_core/SB2/n1769 ), .Y(\U1/aes_core/SB2/n3281 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1413  ( .A(\U1/aes_core/SB2/n3281 ), .Y(
        \U1/aes_core/SB2/n3331 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U1412  ( .A0(\U1/aes_core/SB2/n1976 ), 
        .A1(\U1/aes_core/SB2/n2068 ), .B0(\U1/aes_core/SB2/n3340 ), .B1(
        \U1/aes_core/SB2/n2055 ), .C0(\U1/aes_core/SB2/n3331 ), .C1(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n1777 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1411  ( .A(\U1/aes_core/SB2/n3300 ), .Y(
        \U1/aes_core/SB2/n1952 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1410  ( .A(\U1/aes_core/SB2/n1774 ), .B(
        \U1/aes_core/SB2/n1781 ), .Y(\U1/aes_core/SB2/n2070 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1409  ( .A(\U1/aes_core/SB2/n1770 ), .B(
        \U1/aes_core/SB2/n1769 ), .Y(\U1/aes_core/SB2/n3279 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1408  ( .A0(\U1/aes_core/SB2/n2070 ), 
        .A1(\U1/aes_core/SB2/n3346 ), .B0(\U1/aes_core/SB2/n3279 ), .B1(
        \U1/aes_core/SB2/n1995 ), .Y(\U1/aes_core/SB2/n1771 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1407  ( .A0(\U1/aes_core/SB2/n2058 ), 
        .A1(\U1/aes_core/SB2/n3305 ), .B0(\U1/aes_core/SB2/n1952 ), .B1(
        \U1/aes_core/SB2/n2019 ), .C0(\U1/aes_core/SB2/n1771 ), .Y(
        \U1/aes_core/SB2/n1776 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1406  ( .A(\U1/aes_core/SB2/n3268 ), .B(
        \U1/aes_core/SB2/n2019 ), .Y(\U1/aes_core/SB2/n1880 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1405  ( .A(\U1/aes_core/SB2/n1773 ), .B(
        \U1/aes_core/SB2/n1772 ), .Y(\U1/aes_core/SB2/n3302 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1404  ( .A(\U1/aes_core/SB2/n3302 ), .Y(
        \U1/aes_core/SB2/n3276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1403  ( .A(\U1/aes_core/SB2/n3276 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n1845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1402  ( .A(\U1/aes_core/SB2/n2070 ), .Y(
        \U1/aes_core/SB2/n3324 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1401  ( .A(\U1/aes_core/SB2/n3324 ), .B(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n1929 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1400  ( .A(\U1/aes_core/SB2/n1783 ), .B(
        \U1/aes_core/SB2/n1774 ), .Y(\U1/aes_core/SB2/n2065 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1399  ( .A(\U1/aes_core/SB2/n2065 ), .Y(
        \U1/aes_core/SB2/n3322 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1398  ( .A(\U1/aes_core/SB2/n3322 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1852 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB2/U1397  ( .A(\U1/aes_core/SB2/n1880 ), .B(
        \U1/aes_core/SB2/n1845 ), .C(\U1/aes_core/SB2/n1929 ), .D(
        \U1/aes_core/SB2/n1852 ), .Y(\U1/aes_core/SB2/n1775 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1396  ( .AN(\U1/aes_core/SB2/n1778 ), 
        .B(\U1/aes_core/SB2/n1777 ), .C(\U1/aes_core/SB2/n1776 ), .D(
        \U1/aes_core/SB2/n1775 ), .Y(\U1/aes_core/SB2/n3295 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1395  ( .A(\U1/aes_core/SB2/n1780 ), .B(
        \U1/aes_core/SB2/n1779 ), .Y(\U1/aes_core/SB2/n3297 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1394  ( .A(\U1/aes_core/SB2/n3297 ), .B(
        \U1/aes_core/SB2/n2021 ), .Y(\U1/aes_core/SB2/n1965 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1393  ( .A(\U1/aes_core/SB2/n3300 ), .B(
        \U1/aes_core/SB2/n2006 ), .Y(\U1/aes_core/SB2/n1878 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1392  ( .A(\U1/aes_core/SB2/n3333 ), .B(
        \U1/aes_core/SB2/n3305 ), .Y(\U1/aes_core/SB2/n1842 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1391  ( .A0(\U1/aes_core/SB2/n3300 ), 
        .A1(\U1/aes_core/SB2/n3342 ), .B0(\U1/aes_core/SB2/n1842 ), .Y(
        \U1/aes_core/SB2/n1787 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1390  ( .A(\U1/aes_core/SB2/n1912 ), .Y(
        \U1/aes_core/SB2/n3325 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1389  ( .A(\U1/aes_core/SB2/n3268 ), .B(
        \U1/aes_core/SB2/n3325 ), .Y(\U1/aes_core/SB2/n1977 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1388  ( .A(\U1/aes_core/SB2/n3268 ), .B(
        \U1/aes_core/SB2/n3334 ), .Y(\U1/aes_core/SB2/n1954 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1387  ( .A(\U1/aes_core/SB2/n1782 ), .B(
        \U1/aes_core/SB2/n1781 ), .Y(\U1/aes_core/SB2/n2008 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1386  ( .A(\U1/aes_core/SB2/n2008 ), .Y(
        \U1/aes_core/SB2/n3307 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1385  ( .A(\U1/aes_core/SB2/n3307 ), .B(
        \U1/aes_core/SB2/n2019 ), .Y(\U1/aes_core/SB2/n1855 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1384  ( .A(\U1/aes_core/SB2/n3307 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1902 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1383  ( .A(\U1/aes_core/SB2/n1977 ), .B(
        \U1/aes_core/SB2/n1954 ), .C(\U1/aes_core/SB2/n1855 ), .D(
        \U1/aes_core/SB2/n1902 ), .Y(\U1/aes_core/SB2/n1786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1382  ( .A(\U1/aes_core/SB2/n3346 ), .Y(
        \U1/aes_core/SB2/n3275 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1381  ( .A(\U1/aes_core/SB2/n3275 ), .B(
        \U1/aes_core/SB2/n1976 ), .Y(\U1/aes_core/SB2/n1927 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1380  ( .A(\U1/aes_core/SB2/n3297 ), .Y(
        \U1/aes_core/SB2/n3282 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1379  ( .A(\U1/aes_core/SB2/n1976 ), .B(
        \U1/aes_core/SB2/n3282 ), .Y(\U1/aes_core/SB2/n1922 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1378  ( .A(\U1/aes_core/SB2/n3322 ), .B(
        \U1/aes_core/SB2/n3276 ), .Y(\U1/aes_core/SB2/n1830 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1377  ( .A(\U1/aes_core/SB2/n3299 ), .B(
        \U1/aes_core/SB2/n2019 ), .Y(\U1/aes_core/SB2/n1909 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1376  ( .A(\U1/aes_core/SB2/n1927 ), .B(
        \U1/aes_core/SB2/n1922 ), .C(\U1/aes_core/SB2/n1830 ), .D(
        \U1/aes_core/SB2/n1909 ), .Y(\U1/aes_core/SB2/n1785 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1375  ( .A(\U1/aes_core/SB2/n3279 ), .Y(
        \U1/aes_core/SB2/n3323 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1374  ( .A(\U1/aes_core/SB2/n3274 ), .B(
        \U1/aes_core/SB2/n3323 ), .Y(\U1/aes_core/SB2/n1820 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1373  ( .A(\U1/aes_core/SB2/n2054 ), .B(
        \U1/aes_core/SB2/n3274 ), .Y(\U1/aes_core/SB2/n1864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1372  ( .A(\U1/aes_core/SB2/n1783 ), .B(
        \U1/aes_core/SB2/n1782 ), .Y(\U1/aes_core/SB2/n3303 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1371  ( .A(\U1/aes_core/SB2/n3303 ), .Y(
        \U1/aes_core/SB2/n3329 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1370  ( .A(\U1/aes_core/SB2/n2068 ), .B(
        \U1/aes_core/SB2/n3329 ), .Y(\U1/aes_core/SB2/n1890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1369  ( .A(\U1/aes_core/SB2/n2054 ), .B(
        \U1/aes_core/SB2/n3324 ), .Y(\U1/aes_core/SB2/n1990 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1368  ( .A(\U1/aes_core/SB2/n1820 ), .B(
        \U1/aes_core/SB2/n1864 ), .C(\U1/aes_core/SB2/n1890 ), .D(
        \U1/aes_core/SB2/n1990 ), .Y(\U1/aes_core/SB2/n1784 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1367  ( .A(\U1/aes_core/SB2/n1965 ), .B(
        \U1/aes_core/SB2/n1878 ), .C(\U1/aes_core/SB2/n1787 ), .D(
        \U1/aes_core/SB2/n1786 ), .E(\U1/aes_core/SB2/n1785 ), .F(
        \U1/aes_core/SB2/n1784 ), .Y(\U1/aes_core/SB2/n3286 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1366  ( .A(\U1/aes_core/SB2/n3279 ), .B(
        \U1/aes_core/SB2/n2021 ), .Y(\U1/aes_core/SB2/n1831 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1365  ( .A(\U1/aes_core/SB2/n3280 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n1980 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1364  ( .A(\U1/aes_core/SB2/n3278 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n1872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1363  ( .A(\U1/aes_core/SB2/n3278 ), .B(
        \U1/aes_core/SB2/n3281 ), .Y(\U1/aes_core/SB2/n1881 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1362  ( .A(\U1/aes_core/SB2/n3342 ), .B(
        \U1/aes_core/SB2/n3308 ), .Y(\U1/aes_core/SB2/n1919 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1361  ( .A(\U1/aes_core/SB2/n3307 ), .B(
        \U1/aes_core/SB2/n3325 ), .Y(\U1/aes_core/SB2/n1923 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1360  ( .A(\U1/aes_core/SB2/n2058 ), .B(
        \U1/aes_core/SB2/n3329 ), .Y(\U1/aes_core/SB2/n1844 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1359  ( .A(\U1/aes_core/SB2/n3331 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1857 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1358  ( .AN(\U1/aes_core/SB2/n1919 ), 
        .B(\U1/aes_core/SB2/n1923 ), .C(\U1/aes_core/SB2/n1844 ), .D(
        \U1/aes_core/SB2/n1857 ), .Y(\U1/aes_core/SB2/n1791 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1357  ( .A(\U1/aes_core/SB2/n3300 ), .B(
        \U1/aes_core/SB2/n3281 ), .Y(\U1/aes_core/SB2/n1891 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1356  ( .A(\U1/aes_core/SB2/n3347 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n1967 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1355  ( .A(\U1/aes_core/SB2/n1995 ), .B(
        \U1/aes_core/SB2/n3346 ), .Y(\U1/aes_core/SB2/n1930 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1354  ( .A(\U1/aes_core/SB2/n1995 ), .B(
        \U1/aes_core/SB2/n2006 ), .Y(\U1/aes_core/SB2/n1828 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1353  ( .A0(\U1/aes_core/SB2/n3281 ), 
        .A1(\U1/aes_core/SB2/n1995 ), .B0(\U1/aes_core/SB2/n3300 ), .B1(
        \U1/aes_core/SB2/n3346 ), .Y(\U1/aes_core/SB2/n1789 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1352  ( .A0(\U1/aes_core/SB2/n1888 ), 
        .A1(\U1/aes_core/SB2/n2070 ), .B0(\U1/aes_core/SB2/n2020 ), .B1(
        \U1/aes_core/SB2/n3280 ), .Y(\U1/aes_core/SB2/n1788 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1351  ( .A(\U1/aes_core/SB2/n1891 ), .B(
        \U1/aes_core/SB2/n1967 ), .C(\U1/aes_core/SB2/n1930 ), .D(
        \U1/aes_core/SB2/n1828 ), .E(\U1/aes_core/SB2/n1789 ), .F(
        \U1/aes_core/SB2/n1788 ), .Y(\U1/aes_core/SB2/n1790 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1350  ( .A(\U1/aes_core/SB2/n1831 ), .B(
        \U1/aes_core/SB2/n1980 ), .C(\U1/aes_core/SB2/n1872 ), .D(
        \U1/aes_core/SB2/n1881 ), .E(\U1/aes_core/SB2/n1791 ), .F(
        \U1/aes_core/SB2/n1790 ), .Y(\U1/aes_core/SB2/n3321 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U1349  ( .A1N(\U1/aes_core/SB2/n3299 ), 
        .A0(\U1/aes_core/SB2/n3343 ), .B0(\U1/aes_core/SB2/n2020 ), .Y(
        \U1/aes_core/SB2/n1792 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1348  ( .A(\U1/aes_core/SB2/n1995 ), .B(
        \U1/aes_core/SB2/n2039 ), .Y(\U1/aes_core/SB2/n1943 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1347  ( .A(\U1/aes_core/SB2/n3280 ), .B(
        \U1/aes_core/SB2/n2057 ), .Y(\U1/aes_core/SB2/n1850 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1346  ( .A(\U1/aes_core/SB2/n3280 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n1886 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1345  ( .A(\U1/aes_core/SB2/n1792 ), .B(
        \U1/aes_core/SB2/n1943 ), .C(\U1/aes_core/SB2/n1850 ), .D(
        \U1/aes_core/SB2/n1886 ), .Y(\U1/aes_core/SB2/n1797 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1344  ( .A0(\U1/aes_core/SB2/n2057 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n2021 ), .B1(
        \U1/aes_core/SB2/n3296 ), .C0(\U1/aes_core/SB2/n1912 ), .C1(
        \U1/aes_core/SB2/n3309 ), .Y(\U1/aes_core/SB2/n1796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1343  ( .A(\U1/aes_core/SB2/n3342 ), .B(
        \U1/aes_core/SB2/n3309 ), .Y(\U1/aes_core/SB2/n1972 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1342  ( .A(\U1/aes_core/SB2/n2065 ), .B(
        \U1/aes_core/SB2/n2010 ), .Y(\U1/aes_core/SB2/n1833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1341  ( .A(\U1/aes_core/SB2/n1833 ), .Y(
        \U1/aes_core/SB2/n1793 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1340  ( .A(\U1/aes_core/SB2/n3329 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1339  ( .A(\U1/aes_core/SB2/n1976 ), .B(
        \U1/aes_core/SB2/n2054 ), .Y(\U1/aes_core/SB2/n1853 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1338  ( .AN(\U1/aes_core/SB2/n1972 ), 
        .B(\U1/aes_core/SB2/n1793 ), .C(\U1/aes_core/SB2/n1866 ), .D(
        \U1/aes_core/SB2/n1853 ), .Y(\U1/aes_core/SB2/n1795 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1337  ( .A(\U1/aes_core/SB2/n1888 ), .B(
        \U1/aes_core/SB2/n2021 ), .Y(\U1/aes_core/SB2/n1918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1336  ( .A(\U1/aes_core/SB2/n1806 ), .B(
        \U1/aes_core/SB2/n3297 ), .Y(\U1/aes_core/SB2/n1895 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1335  ( .A(\U1/aes_core/SB2/n2008 ), .B(
        \U1/aes_core/SB2/n2020 ), .Y(\U1/aes_core/SB2/n1935 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1334  ( .A(\U1/aes_core/SB2/n2008 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n1827 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1333  ( .A(\U1/aes_core/SB2/n1918 ), .B(
        \U1/aes_core/SB2/n1895 ), .C(\U1/aes_core/SB2/n1935 ), .D(
        \U1/aes_core/SB2/n1827 ), .Y(\U1/aes_core/SB2/n1794 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1332  ( .A(\U1/aes_core/SB2/n1797 ), .B(
        \U1/aes_core/SB2/n1796 ), .C(\U1/aes_core/SB2/n1795 ), .D(
        \U1/aes_core/SB2/n1794 ), .Y(\U1/aes_core/SB2/n3293 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1331  ( .A(\U1/aes_core/SB2/n3308 ), .Y(
        \U1/aes_core/SB2/n3327 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1330  ( .A0(\U1/aes_core/SB2/n3330 ), 
        .A1(\U1/aes_core/SB2/n3268 ), .B0(\U1/aes_core/SB2/n2068 ), .B1(
        \U1/aes_core/SB2/n3327 ), .Y(\U1/aes_core/SB2/n1798 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1329  ( .A0(\U1/aes_core/SB2/n3297 ), 
        .A1(\U1/aes_core/SB2/n3347 ), .B0(\U1/aes_core/SB2/n3280 ), .B1(
        \U1/aes_core/SB2/n3346 ), .C0(\U1/aes_core/SB2/n1798 ), .Y(
        \U1/aes_core/SB2/n1804 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1328  ( .A(\U1/aes_core/SB2/n3303 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n1862 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1327  ( .A(\U1/aes_core/SB2/n3332 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1326  ( .A(\U1/aes_core/SB2/n3268 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1325  ( .A(\U1/aes_core/SB2/n3330 ), .B(
        \U1/aes_core/SB2/n3307 ), .Y(\U1/aes_core/SB2/n1839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1324  ( .AN(\U1/aes_core/SB2/n1862 ), 
        .B(\U1/aes_core/SB2/n1874 ), .C(\U1/aes_core/SB2/n1867 ), .D(
        \U1/aes_core/SB2/n1839 ), .Y(\U1/aes_core/SB2/n1803 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1323  ( .A(\U1/aes_core/SB2/n3281 ), .B(
        \U1/aes_core/SB2/n2057 ), .Y(\U1/aes_core/SB2/n1948 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1322  ( .A0(\U1/aes_core/SB2/n3325 ), 
        .A1(\U1/aes_core/SB2/n1948 ), .B0(\U1/aes_core/SB2/n3322 ), .Y(
        \U1/aes_core/SB2/n1801 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1321  ( .A(\U1/aes_core/SB2/n3344 ), .Y(
        \U1/aes_core/SB2/n1949 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1320  ( .A0(\U1/aes_core/SB2/n2058 ), 
        .A1(\U1/aes_core/SB2/n3323 ), .B0(\U1/aes_core/SB2/n1949 ), .Y(
        \U1/aes_core/SB2/n1800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1319  ( .A(\U1/aes_core/SB2/n2020 ), .Y(
        \U1/aes_core/SB2/n2060 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1318  ( .A0(\U1/aes_core/SB2/n1952 ), 
        .A1(\U1/aes_core/SB2/n1976 ), .B0(\U1/aes_core/SB2/n2060 ), .Y(
        \U1/aes_core/SB2/n1799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1317  ( .A(\U1/aes_core/SB2/n2058 ), .B(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n1925 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1316  ( .A(\U1/aes_core/SB2/n1801 ), .B(
        \U1/aes_core/SB2/n1800 ), .C(\U1/aes_core/SB2/n1799 ), .D(
        \U1/aes_core/SB2/n1925 ), .Y(\U1/aes_core/SB2/n1802 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1315  ( .A(\U1/aes_core/SB2/n3286 ), .B(
        \U1/aes_core/SB2/n3321 ), .C(\U1/aes_core/SB2/n3293 ), .D(
        \U1/aes_core/SB2/n1804 ), .E(\U1/aes_core/SB2/n1803 ), .F(
        \U1/aes_core/SB2/n1802 ), .Y(\U1/aes_core/SB2/n2074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1314  ( .A0(\U1/aes_core/SB2/n2019 ), 
        .A1(\U1/aes_core/SB2/n3330 ), .B0(\U1/aes_core/SB2/n3324 ), .Y(
        \U1/aes_core/SB2/n1805 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1313  ( .A(\U1/aes_core/SB2/n3269 ), .B(
        \U1/aes_core/SB2/n2058 ), .Y(\U1/aes_core/SB2/n1910 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1312  ( .A(\U1/aes_core/SB2/n2055 ), .B(
        \U1/aes_core/SB2/n3276 ), .Y(\U1/aes_core/SB2/n1819 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1311  ( .A(\U1/aes_core/SB2/n3340 ), .B(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n1921 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1310  ( .A(\U1/aes_core/SB2/n1805 ), .B(
        \U1/aes_core/SB2/n1910 ), .C(\U1/aes_core/SB2/n1819 ), .D(
        \U1/aes_core/SB2/n1921 ), .Y(\U1/aes_core/SB2/n1810 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1309  ( .A0(\U1/aes_core/SB2/n2020 ), 
        .A1(\U1/aes_core/SB2/n1806 ), .B0(\U1/aes_core/SB2/n3302 ), .B1(
        \U1/aes_core/SB2/n3347 ), .C0(\U1/aes_core/SB2/n3346 ), .C1(
        \U1/aes_core/SB2/n2065 ), .Y(\U1/aes_core/SB2/n1809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1308  ( .A(\U1/aes_core/SB2/n1976 ), .B(
        \U1/aes_core/SB2/n3334 ), .Y(\U1/aes_core/SB2/n1841 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1307  ( .A(\U1/aes_core/SB2/n2058 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1964 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1306  ( .A(\U1/aes_core/SB2/n3275 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1863 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1305  ( .A(\U1/aes_core/SB2/n3340 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1926 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1304  ( .A(\U1/aes_core/SB2/n1841 ), .B(
        \U1/aes_core/SB2/n1964 ), .C(\U1/aes_core/SB2/n1863 ), .D(
        \U1/aes_core/SB2/n1926 ), .Y(\U1/aes_core/SB2/n1808 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1303  ( .A(\U1/aes_core/SB2/n3340 ), .B(
        \U1/aes_core/SB2/n3332 ), .Y(\U1/aes_core/SB2/n1889 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1302  ( .A(\U1/aes_core/SB2/n3333 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n1876 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1301  ( .A(\U1/aes_core/SB2/n3274 ), .B(
        \U1/aes_core/SB2/n3276 ), .Y(\U1/aes_core/SB2/n1854 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1300  ( .A(\U1/aes_core/SB2/n3323 ), .B(
        \U1/aes_core/SB2/n3327 ), .Y(\U1/aes_core/SB2/n1829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1299  ( .A(\U1/aes_core/SB2/n1889 ), .B(
        \U1/aes_core/SB2/n1876 ), .C(\U1/aes_core/SB2/n1854 ), .D(
        \U1/aes_core/SB2/n1829 ), .Y(\U1/aes_core/SB2/n1807 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1298  ( .A(\U1/aes_core/SB2/n1810 ), .B(
        \U1/aes_core/SB2/n1809 ), .C(\U1/aes_core/SB2/n1808 ), .D(
        \U1/aes_core/SB2/n1807 ), .Y(\U1/aes_core/SB2/n1811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1297  ( .A(\U1/aes_core/SB2/n1811 ), .Y(
        \U1/aes_core/SB2/n3284 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1296  ( .A0(\U1/aes_core/SB2/n3308 ), 
        .A1(\U1/aes_core/SB2/n2039 ), .B0(\U1/aes_core/SB2/n3297 ), .B1(
        \U1/aes_core/SB2/n2070 ), .C0(\U1/aes_core/SB2/n3284 ), .Y(
        \U1/aes_core/SB2/n1818 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1295  ( .A(\U1/aes_core/SB2/n3329 ), .B(
        \U1/aes_core/SB2/n3274 ), .Y(\U1/aes_core/SB2/n1920 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U1294  ( .A1N(\U1/aes_core/SB2/n1920 ), 
        .A0(\U1/aes_core/SB2/n3305 ), .B0(\U1/aes_core/SB2/n2019 ), .Y(
        \U1/aes_core/SB2/n1814 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1293  ( .A(\U1/aes_core/SB2/n2017 ), .B(
        \U1/aes_core/SB2/n3346 ), .Y(\U1/aes_core/SB2/n2018 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1292  ( .A0(\U1/aes_core/SB2/n3331 ), 
        .A1(\U1/aes_core/SB2/n2018 ), .B0(\U1/aes_core/SB2/n3268 ), .Y(
        \U1/aes_core/SB2/n1813 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1291  ( .A0(\U1/aes_core/SB2/n2058 ), 
        .A1(\U1/aes_core/SB2/n3333 ), .B0(\U1/aes_core/SB2/n2055 ), .Y(
        \U1/aes_core/SB2/n1812 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1290  ( .A(\U1/aes_core/SB2/n2054 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n1851 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1289  ( .A(\U1/aes_core/SB2/n1814 ), .B(
        \U1/aes_core/SB2/n1813 ), .C(\U1/aes_core/SB2/n1812 ), .D(
        \U1/aes_core/SB2/n1851 ), .Y(\U1/aes_core/SB2/n1817 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1288  ( .A(\U1/aes_core/SB2/n3275 ), .B(
        \U1/aes_core/SB2/n2060 ), .Y(\U1/aes_core/SB2/n2059 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1287  ( .A(\U1/aes_core/SB2/n2053 ), .B(
        \U1/aes_core/SB2/n1976 ), .Y(\U1/aes_core/SB2/n1815 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1286  ( .A0(\U1/aes_core/SB2/n2059 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n1815 ), .B1(
        \U1/aes_core/SB2/n2010 ), .C0(\U1/aes_core/SB2/n3302 ), .C1(
        \U1/aes_core/SB2/n3278 ), .Y(\U1/aes_core/SB2/n1816 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1285  ( .A(\U1/aes_core/SB2/n3353 ), .B(
        \U1/aes_core/SB2/n3295 ), .C(\U1/aes_core/SB2/n2074 ), .D(
        \U1/aes_core/SB2/n1818 ), .E(\U1/aes_core/SB2/n1817 ), .F(
        \U1/aes_core/SB2/n1816 ), .Y(\U1/aes_core/sb2 [10]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1284  ( .A(\U1/aes_core/SB2/n3347 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n2034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1283  ( .A(\U1/aes_core/SB2/n3330 ), .B(
        \U1/aes_core/SB2/n1952 ), .Y(\U1/aes_core/SB2/n2036 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1282  ( .AN(\U1/aes_core/SB2/n1821 ), 
        .B(\U1/aes_core/SB2/n1820 ), .C(\U1/aes_core/SB2/n1819 ), .D(
        \U1/aes_core/SB2/n2036 ), .Y(\U1/aes_core/SB2/n1826 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1281  ( .A(\U1/aes_core/SB2/n3324 ), .B(
        \U1/aes_core/SB2/n2055 ), .Y(\U1/aes_core/SB2/n1983 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1280  ( .A0(\U1/aes_core/SB2/n3269 ), 
        .A1(\U1/aes_core/SB2/n3268 ), .B0(\U1/aes_core/SB2/n3323 ), .Y(
        \U1/aes_core/SB2/n1822 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1279  ( .A(\U1/aes_core/SB2/n3340 ), .B(
        \U1/aes_core/SB2/n1952 ), .Y(\U1/aes_core/SB2/n2061 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U1278  ( .A0(\U1/aes_core/SB2/n1983 ), 
        .A1(\U1/aes_core/SB2/n3296 ), .B0(\U1/aes_core/SB2/n1822 ), .C0(
        \U1/aes_core/SB2/n2061 ), .Y(\U1/aes_core/SB2/n1825 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1277  ( .A0(\U1/aes_core/SB2/n2020 ), 
        .A1(\U1/aes_core/SB2/n2070 ), .B0(\U1/aes_core/SB2/n1823 ), .B1(
        \U1/aes_core/SB2/n3308 ), .C0(\U1/aes_core/SB2/n3281 ), .C1(
        \U1/aes_core/SB2/n2065 ), .Y(\U1/aes_core/SB2/n1824 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1276  ( .A(\U1/aes_core/SB2/n1828 ), .B(
        \U1/aes_core/SB2/n2034 ), .C(\U1/aes_core/SB2/n1827 ), .D(
        \U1/aes_core/SB2/n1826 ), .E(\U1/aes_core/SB2/n1825 ), .F(
        \U1/aes_core/SB2/n1824 ), .Y(\U1/aes_core/SB2/n1962 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1275  ( .A(\U1/aes_core/SB2/n3323 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n2040 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1274  ( .AN(\U1/aes_core/SB2/n1831 ), 
        .B(\U1/aes_core/SB2/n1830 ), .C(\U1/aes_core/SB2/n1829 ), .D(
        \U1/aes_core/SB2/n2040 ), .Y(\U1/aes_core/SB2/n1838 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U1273  ( .A0(\U1/aes_core/SB2/n3331 ), 
        .A1(\U1/aes_core/SB2/n3327 ), .B0(\U1/aes_core/SB2/n3332 ), .B1(
        \U1/aes_core/SB2/n3334 ), .C0(\U1/aes_core/SB2/n3274 ), .C1(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n1837 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1272  ( .A0(\U1/aes_core/SB2/n3301 ), 
        .A1(\U1/aes_core/SB2/n3280 ), .B0(\U1/aes_core/SB2/n2021 ), .B1(
        \U1/aes_core/SB2/n2020 ), .Y(\U1/aes_core/SB2/n1832 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1271  ( .A0(\U1/aes_core/SB2/n1952 ), 
        .A1(\U1/aes_core/SB2/n3323 ), .B0(\U1/aes_core/SB2/n3276 ), .B1(
        \U1/aes_core/SB2/n3299 ), .C0(\U1/aes_core/SB2/n1832 ), .Y(
        \U1/aes_core/SB2/n1836 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1270  ( .A(\U1/aes_core/SB2/n3308 ), .B(
        \U1/aes_core/SB2/n3343 ), .Y(\U1/aes_core/SB2/n3270 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1269  ( .A(\U1/aes_core/SB2/n3344 ), .B(
        \U1/aes_core/SB2/n3347 ), .Y(\U1/aes_core/SB2/n1834 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1268  ( .A0(\U1/aes_core/SB2/n3340 ), 
        .A1(\U1/aes_core/SB2/n3270 ), .B0(\U1/aes_core/SB2/n2058 ), .B1(
        \U1/aes_core/SB2/n1834 ), .C0(\U1/aes_core/SB2/n1833 ), .Y(
        \U1/aes_core/SB2/n1835 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1267  ( .AN(\U1/aes_core/SB2/n1838 ), 
        .B(\U1/aes_core/SB2/n1837 ), .C(\U1/aes_core/SB2/n1836 ), .D(
        \U1/aes_core/SB2/n1835 ), .Y(\U1/aes_core/SB2/n1988 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1266  ( .A(\U1/aes_core/SB2/n1995 ), .B(
        \U1/aes_core/SB2/n3302 ), .Y(\U1/aes_core/SB2/n2024 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1265  ( .A0(\U1/aes_core/SB2/n3303 ), 
        .A1(\U1/aes_core/SB2/n3302 ), .B0(\U1/aes_core/SB2/n1839 ), .Y(
        \U1/aes_core/SB2/n1849 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1264  ( .A0(\U1/aes_core/SB2/n2058 ), 
        .A1(\U1/aes_core/SB2/n3332 ), .B0(\U1/aes_core/SB2/n3275 ), .B1(
        \U1/aes_core/SB2/n3307 ), .Y(\U1/aes_core/SB2/n1840 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1263  ( .A0(\U1/aes_core/SB2/n3344 ), 
        .A1(\U1/aes_core/SB2/n2039 ), .B0(\U1/aes_core/SB2/n2057 ), .B1(
        \U1/aes_core/SB2/n3343 ), .C0(\U1/aes_core/SB2/n1840 ), .Y(
        \U1/aes_core/SB2/n1848 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1262  ( .A(\U1/aes_core/SB2/n1912 ), .B(
        \U1/aes_core/SB2/n3308 ), .Y(\U1/aes_core/SB2/n3292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1261  ( .A(\U1/aes_core/SB2/n3305 ), .B(
        \U1/aes_core/SB2/n3323 ), .Y(\U1/aes_core/SB2/n2037 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1260  ( .AN(\U1/aes_core/SB2/n3292 ), 
        .B(\U1/aes_core/SB2/n1842 ), .C(\U1/aes_core/SB2/n1841 ), .D(
        \U1/aes_core/SB2/n2037 ), .Y(\U1/aes_core/SB2/n1847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1259  ( .A(\U1/aes_core/SB2/n3280 ), .B(
        \U1/aes_core/SB2/n3297 ), .Y(\U1/aes_core/SB2/n2015 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1258  ( .AN(\U1/aes_core/SB2/n2015 ), 
        .B(\U1/aes_core/SB2/n1845 ), .C(\U1/aes_core/SB2/n1844 ), .D(
        \U1/aes_core/SB2/n1843 ), .Y(\U1/aes_core/SB2/n1846 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1257  ( .A(\U1/aes_core/SB2/n2024 ), .B(
        \U1/aes_core/SB2/n1850 ), .C(\U1/aes_core/SB2/n1849 ), .D(
        \U1/aes_core/SB2/n1848 ), .E(\U1/aes_core/SB2/n1847 ), .F(
        \U1/aes_core/SB2/n1846 ), .Y(\U1/aes_core/SB2/n1924 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1256  ( .A(\U1/aes_core/SB2/n2017 ), .B(
        \U1/aes_core/SB2/n3300 ), .Y(\U1/aes_core/SB2/n2064 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1255  ( .A0(\U1/aes_core/SB2/n2017 ), 
        .A1(\U1/aes_core/SB2/n3280 ), .B0(\U1/aes_core/SB2/n1851 ), .Y(
        \U1/aes_core/SB2/n1861 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1254  ( .A(\U1/aes_core/SB2/n3343 ), .B(
        \U1/aes_core/SB2/n1912 ), .Y(\U1/aes_core/SB2/n2023 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1253  ( .A(\U1/aes_core/SB2/n1949 ), .B(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n3312 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1252  ( .AN(\U1/aes_core/SB2/n2023 ), 
        .B(\U1/aes_core/SB2/n1853 ), .C(\U1/aes_core/SB2/n1852 ), .D(
        \U1/aes_core/SB2/n3312 ), .Y(\U1/aes_core/SB2/n1860 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1251  ( .A(\U1/aes_core/SB2/n3274 ), .B(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n2045 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1250  ( .A(\U1/aes_core/SB2/n3339 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n3267 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1249  ( .A(\U1/aes_core/SB2/n2019 ), .B(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n3335 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1248  ( .A(\U1/aes_core/SB2/n1854 ), .B(
        \U1/aes_core/SB2/n2045 ), .C(\U1/aes_core/SB2/n3267 ), .D(
        \U1/aes_core/SB2/n3335 ), .Y(\U1/aes_core/SB2/n1859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1247  ( .A(\U1/aes_core/SB2/n3322 ), .B(
        \U1/aes_core/SB2/n3333 ), .Y(\U1/aes_core/SB2/n2005 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1246  ( .A(\U1/aes_core/SB2/n1857 ), .B(
        \U1/aes_core/SB2/n1856 ), .C(\U1/aes_core/SB2/n2005 ), .D(
        \U1/aes_core/SB2/n1855 ), .Y(\U1/aes_core/SB2/n1858 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1245  ( .A(\U1/aes_core/SB2/n2064 ), .B(
        \U1/aes_core/SB2/n1862 ), .C(\U1/aes_core/SB2/n1861 ), .D(
        \U1/aes_core/SB2/n1860 ), .E(\U1/aes_core/SB2/n1859 ), .F(
        \U1/aes_core/SB2/n1858 ), .Y(\U1/aes_core/SB2/n1940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1244  ( .A(\U1/aes_core/SB2/n3302 ), .B(
        \U1/aes_core/SB2/n2021 ), .Y(\U1/aes_core/SB2/n2016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1243  ( .A(\U1/aes_core/SB2/n3324 ), .B(
        \U1/aes_core/SB2/n3331 ), .Y(\U1/aes_core/SB2/n2041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1242  ( .A(\U1/aes_core/SB2/n3334 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n3265 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1241  ( .A(\U1/aes_core/SB2/n1864 ), .B(
        \U1/aes_core/SB2/n1863 ), .C(\U1/aes_core/SB2/n2041 ), .D(
        \U1/aes_core/SB2/n3265 ), .Y(\U1/aes_core/SB2/n1871 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1240  ( .A(\U1/aes_core/SB2/n1952 ), .B(
        \U1/aes_core/SB2/n3276 ), .Y(\U1/aes_core/SB2/n2027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1239  ( .A(\U1/aes_core/SB2/n3333 ), .B(
        \U1/aes_core/SB2/n1952 ), .Y(\U1/aes_core/SB2/n3311 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1238  ( .A(\U1/aes_core/SB2/n1866 ), .B(
        \U1/aes_core/SB2/n2027 ), .C(\U1/aes_core/SB2/n1865 ), .D(
        \U1/aes_core/SB2/n3311 ), .Y(\U1/aes_core/SB2/n1870 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U1237  ( .A(\U1/aes_core/SB2/n2055 ), .B(
        \U1/aes_core/SB2/n3329 ), .C(\U1/aes_core/SB2/n2053 ), .Y(
        \U1/aes_core/SB2/n1868 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1236  ( .A0(\U1/aes_core/SB2/n1868 ), 
        .A1(\U1/aes_core/SB2/n2010 ), .B0(\U1/aes_core/SB2/n2020 ), .B1(
        \U1/aes_core/SB2/n3347 ), .C0(\U1/aes_core/SB2/n1867 ), .Y(
        \U1/aes_core/SB2/n1869 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1235  ( .A(\U1/aes_core/SB2/n2016 ), .B(
        \U1/aes_core/SB2/n1873 ), .C(\U1/aes_core/SB2/n1872 ), .D(
        \U1/aes_core/SB2/n1871 ), .E(\U1/aes_core/SB2/n1870 ), .F(
        \U1/aes_core/SB2/n1869 ), .Y(\U1/aes_core/SB2/n1973 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1234  ( .A(\U1/aes_core/SB2/n3300 ), .B(
        \U1/aes_core/SB2/n1888 ), .Y(\U1/aes_core/SB2/n2028 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1233  ( .A0(\U1/aes_core/SB2/n2020 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n1874 ), .Y(
        \U1/aes_core/SB2/n1885 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1232  ( .A0(\U1/aes_core/SB2/n1976 ), 
        .A1(\U1/aes_core/SB2/n2019 ), .B0(\U1/aes_core/SB2/n3322 ), .B1(
        \U1/aes_core/SB2/n3334 ), .Y(\U1/aes_core/SB2/n1875 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1231  ( .A0(\U1/aes_core/SB2/n3308 ), 
        .A1(\U1/aes_core/SB2/n3346 ), .B0(\U1/aes_core/SB2/n3303 ), .B1(
        \U1/aes_core/SB2/n3279 ), .C0(\U1/aes_core/SB2/n1875 ), .Y(
        \U1/aes_core/SB2/n1884 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1230  ( .A(\U1/aes_core/SB2/n3303 ), .B(
        \U1/aes_core/SB2/n2020 ), .Y(\U1/aes_core/SB2/n3291 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1229  ( .A(\U1/aes_core/SB2/n3291 ), .Y(
        \U1/aes_core/SB2/n1877 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1228  ( .A(\U1/aes_core/SB2/n3332 ), .B(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n2047 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1227  ( .AN(\U1/aes_core/SB2/n1878 ), 
        .B(\U1/aes_core/SB2/n1877 ), .C(\U1/aes_core/SB2/n1876 ), .D(
        \U1/aes_core/SB2/n2047 ), .Y(\U1/aes_core/SB2/n1883 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1226  ( .A(\U1/aes_core/SB2/n2058 ), .B(
        \U1/aes_core/SB2/n3307 ), .Y(\U1/aes_core/SB2/n2003 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1225  ( .AN(\U1/aes_core/SB2/n1881 ), 
        .B(\U1/aes_core/SB2/n1880 ), .C(\U1/aes_core/SB2/n1879 ), .D(
        \U1/aes_core/SB2/n2003 ), .Y(\U1/aes_core/SB2/n1882 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1224  ( .A(\U1/aes_core/SB2/n2028 ), .B(
        \U1/aes_core/SB2/n1886 ), .C(\U1/aes_core/SB2/n1885 ), .D(
        \U1/aes_core/SB2/n1884 ), .E(\U1/aes_core/SB2/n1883 ), .F(
        \U1/aes_core/SB2/n1882 ), .Y(\U1/aes_core/SB2/n1947 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1223  ( .A0(\U1/aes_core/SB2/n2053 ), 
        .A1(\U1/aes_core/SB2/n2018 ), .B0(\U1/aes_core/SB2/n1976 ), .B1(
        \U1/aes_core/SB2/n2060 ), .Y(\U1/aes_core/SB2/n1887 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1222  ( .A0(\U1/aes_core/SB2/n3281 ), 
        .A1(\U1/aes_core/SB2/n3280 ), .B0(\U1/aes_core/SB2/n1888 ), .B1(
        \U1/aes_core/SB2/n3343 ), .C0(\U1/aes_core/SB2/n1887 ), .Y(
        \U1/aes_core/SB2/n1898 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1221  ( .A(\U1/aes_core/SB2/n3329 ), .B(
        \U1/aes_core/SB2/n3325 ), .Y(\U1/aes_core/SB2/n2044 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1220  ( .AN(\U1/aes_core/SB2/n1891 ), 
        .B(\U1/aes_core/SB2/n1890 ), .C(\U1/aes_core/SB2/n1889 ), .D(
        \U1/aes_core/SB2/n2044 ), .Y(\U1/aes_core/SB2/n1897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1219  ( .A0(\U1/aes_core/SB2/n3282 ), 
        .A1(\U1/aes_core/SB2/n3340 ), .B0(\U1/aes_core/SB2/n3322 ), .Y(
        \U1/aes_core/SB2/n1894 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1218  ( .A(\U1/aes_core/SB2/n3344 ), .B(
        \U1/aes_core/SB2/n1995 ), .Y(\U1/aes_core/SB2/n1892 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1217  ( .A0(\U1/aes_core/SB2/n3333 ), 
        .A1(\U1/aes_core/SB2/n1892 ), .B0(\U1/aes_core/SB2/n3329 ), .B1(
        \U1/aes_core/SB2/n1948 ), .Y(\U1/aes_core/SB2/n1893 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1216  ( .AN(\U1/aes_core/SB2/n1895 ), 
        .B(\U1/aes_core/SB2/n1894 ), .C(\U1/aes_core/SB2/n1893 ), .Y(
        \U1/aes_core/SB2/n1896 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1215  ( .A(\U1/aes_core/SB2/n1940 ), .B(
        \U1/aes_core/SB2/n1973 ), .C(\U1/aes_core/SB2/n1947 ), .D(
        \U1/aes_core/SB2/n1898 ), .E(\U1/aes_core/SB2/n1897 ), .F(
        \U1/aes_core/SB2/n1896 ), .Y(\U1/aes_core/SB2/n1999 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1214  ( .A(\U1/aes_core/SB2/n1962 ), .B(
        \U1/aes_core/SB2/n1988 ), .C(\U1/aes_core/SB2/n1924 ), .D(
        \U1/aes_core/SB2/n1999 ), .Y(\U1/aes_core/SB2/n1908 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1213  ( .A(\U1/aes_core/SB2/n3333 ), .B(
        \U1/aes_core/SB2/n2068 ), .Y(\U1/aes_core/SB2/n2009 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1212  ( .A(\U1/aes_core/SB2/n3323 ), .B(
        \U1/aes_core/SB2/n2060 ), .Y(\U1/aes_core/SB2/n2002 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1211  ( .A(\U1/aes_core/SB2/n3297 ), .B(
        \U1/aes_core/SB2/n3302 ), .Y(\U1/aes_core/SB2/n3306 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1210  ( .A0(\U1/aes_core/SB2/n1952 ), 
        .A1(\U1/aes_core/SB2/n3275 ), .B0(\U1/aes_core/SB2/n3306 ), .B1(
        \U1/aes_core/SB2/n3305 ), .Y(\U1/aes_core/SB2/n1899 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1209  ( .A0(\U1/aes_core/SB2/n2021 ), 
        .A1(\U1/aes_core/SB2/n2009 ), .B0(\U1/aes_core/SB2/n3278 ), .B1(
        \U1/aes_core/SB2/n2002 ), .C0(\U1/aes_core/SB2/n1899 ), .Y(
        \U1/aes_core/SB2/n1900 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1208  ( .A(\U1/aes_core/SB2/n1900 ), .Y(
        \U1/aes_core/SB2/n1907 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1207  ( .A0(\U1/aes_core/SB2/n3301 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n2020 ), .B1(
        \U1/aes_core/SB2/n1995 ), .Y(\U1/aes_core/SB2/n1901 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1206  ( .A0(\U1/aes_core/SB2/n2054 ), 
        .A1(\U1/aes_core/SB2/n3268 ), .B0(\U1/aes_core/SB2/n3327 ), .B1(
        \U1/aes_core/SB2/n3282 ), .C0(\U1/aes_core/SB2/n1901 ), .Y(
        \U1/aes_core/SB2/n1906 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1205  ( .A0(\U1/aes_core/SB2/n2068 ), 
        .A1(\U1/aes_core/SB2/n3323 ), .B0(\U1/aes_core/SB2/n2055 ), .Y(
        \U1/aes_core/SB2/n1904 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1204  ( .A(\U1/aes_core/SB2/n3340 ), .B(
        \U1/aes_core/SB2/n3305 ), .Y(\U1/aes_core/SB2/n2026 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB2/U1203  ( .A(\U1/aes_core/SB2/n1904 ), .B(
        \U1/aes_core/SB2/n2026 ), .C(\U1/aes_core/SB2/n1903 ), .D(
        \U1/aes_core/SB2/n1902 ), .Y(\U1/aes_core/SB2/n1905 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1202  ( .AN(\U1/aes_core/SB2/n1908 ), 
        .B(\U1/aes_core/SB2/n1907 ), .C(\U1/aes_core/SB2/n1906 ), .D(
        \U1/aes_core/SB2/n1905 ), .Y(\U1/aes_core/sb2 [11]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1201  ( .A0(\U1/aes_core/SB2/n1920 ), 
        .A1(\U1/aes_core/SB2/n2008 ), .B0(\U1/aes_core/SB2/n3297 ), .Y(
        \U1/aes_core/SB2/n1917 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1200  ( .A(\U1/aes_core/SB2/n1949 ), .B(
        \U1/aes_core/SB2/n3325 ), .Y(\U1/aes_core/SB2/n2035 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U1199  ( .A(\U1/aes_core/SB2/n1910 ), .B(
        \U1/aes_core/SB2/n2035 ), .C(\U1/aes_core/SB2/n1909 ), .Y(
        \U1/aes_core/SB2/n1916 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1198  ( .A(\U1/aes_core/SB2/n2053 ), .B(
        \U1/aes_core/SB2/n3322 ), .Y(\U1/aes_core/SB2/n1913 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1197  ( .A(\U1/aes_core/SB2/n3305 ), .B(
        \U1/aes_core/SB2/n1952 ), .Y(\U1/aes_core/SB2/n1911 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1196  ( .A0(\U1/aes_core/SB2/n1913 ), 
        .A1(\U1/aes_core/SB2/n1912 ), .B0(\U1/aes_core/SB2/n1911 ), .B1(
        \U1/aes_core/SB2/n2057 ), .C0(\U1/aes_core/SB2/n2006 ), .C1(
        \U1/aes_core/SB2/n2008 ), .Y(\U1/aes_core/SB2/n1915 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1195  ( .A0(\U1/aes_core/SB2/n3303 ), 
        .A1(\U1/aes_core/SB2/n2017 ), .B0(\U1/aes_core/SB2/n3281 ), .B1(
        \U1/aes_core/SB2/n3343 ), .C0(\U1/aes_core/SB2/n3308 ), .C1(
        \U1/aes_core/SB2/n2010 ), .Y(\U1/aes_core/SB2/n1914 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1194  ( .A(\U1/aes_core/SB2/n1919 ), .B(
        \U1/aes_core/SB2/n1918 ), .C(\U1/aes_core/SB2/n1917 ), .D(
        \U1/aes_core/SB2/n1916 ), .E(\U1/aes_core/SB2/n1915 ), .F(
        \U1/aes_core/SB2/n1914 ), .Y(\U1/aes_core/SB2/n2000 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1193  ( .A0(\U1/aes_core/SB2/n1920 ), 
        .A1(\U1/aes_core/SB2/n3280 ), .B0(\U1/aes_core/SB2/n3346 ), .Y(
        \U1/aes_core/SB2/n1946 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB2/U1192  ( .A0(\U1/aes_core/SB2/n3296 ), 
        .A1(\U1/aes_core/SB2/n3279 ), .A2(\U1/aes_core/SB2/n2010 ), .B0(
        \U1/aes_core/SB2/n3309 ), .Y(\U1/aes_core/SB2/n1945 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1191  ( .A(\U1/aes_core/SB2/n3276 ), .B(
        \U1/aes_core/SB2/n3327 ), .Y(\U1/aes_core/SB2/n2042 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1190  ( .A(\U1/aes_core/SB2/n1923 ), .B(
        \U1/aes_core/SB2/n1922 ), .C(\U1/aes_core/SB2/n1921 ), .D(
        \U1/aes_core/SB2/n2042 ), .Y(\U1/aes_core/SB2/n1942 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1189  ( .A(\U1/aes_core/SB2/n1924 ), .Y(
        \U1/aes_core/SB2/n1939 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1188  ( .A(\U1/aes_core/SB2/n3309 ), .B(
        \U1/aes_core/SB2/n3302 ), .Y(\U1/aes_core/SB2/n2022 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1187  ( .A0(\U1/aes_core/SB2/n2002 ), 
        .A1(\U1/aes_core/SB2/n2065 ), .B0(\U1/aes_core/SB2/n1925 ), .Y(
        \U1/aes_core/SB2/n1934 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1186  ( .A0(\U1/aes_core/SB2/n3280 ), 
        .A1(\U1/aes_core/SB2/n3342 ), .B0(\U1/aes_core/SB2/n3297 ), .B1(
        \U1/aes_core/SB2/n1995 ), .C0(\U1/aes_core/SB2/n3281 ), .C1(
        \U1/aes_core/SB2/n3309 ), .Y(\U1/aes_core/SB2/n1933 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1185  ( .A(\U1/aes_core/SB2/n3307 ), .B(
        \U1/aes_core/SB2/n3323 ), .Y(\U1/aes_core/SB2/n2046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1184  ( .A(\U1/aes_core/SB2/n2068 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n3272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1183  ( .A(\U1/aes_core/SB2/n1927 ), .B(
        \U1/aes_core/SB2/n1926 ), .C(\U1/aes_core/SB2/n2046 ), .D(
        \U1/aes_core/SB2/n3272 ), .Y(\U1/aes_core/SB2/n1932 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1182  ( .A(\U1/aes_core/SB2/n3333 ), .B(
        \U1/aes_core/SB2/n3299 ), .Y(\U1/aes_core/SB2/n2004 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1181  ( .AN(\U1/aes_core/SB2/n1930 ), 
        .B(\U1/aes_core/SB2/n1929 ), .C(\U1/aes_core/SB2/n1928 ), .D(
        \U1/aes_core/SB2/n2004 ), .Y(\U1/aes_core/SB2/n1931 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1180  ( .A(\U1/aes_core/SB2/n2022 ), .B(
        \U1/aes_core/SB2/n1935 ), .C(\U1/aes_core/SB2/n1934 ), .D(
        \U1/aes_core/SB2/n1933 ), .E(\U1/aes_core/SB2/n1932 ), .F(
        \U1/aes_core/SB2/n1931 ), .Y(\U1/aes_core/SB2/n1936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1179  ( .A(\U1/aes_core/SB2/n1936 ), .Y(
        \U1/aes_core/SB2/n1989 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1178  ( .A0(\U1/aes_core/SB2/n3344 ), 
        .A1(\U1/aes_core/SB2/n2017 ), .B0(\U1/aes_core/SB2/n3281 ), .B1(
        \U1/aes_core/SB2/n3347 ), .Y(\U1/aes_core/SB2/n1937 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U1177  ( .A0(\U1/aes_core/SB2/n3324 ), 
        .A1(\U1/aes_core/SB2/n3323 ), .B0(\U1/aes_core/SB2/n3330 ), .B1(
        \U1/aes_core/SB2/n3299 ), .C0(\U1/aes_core/SB2/n1937 ), .Y(
        \U1/aes_core/SB2/n1938 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1176  ( .AN(\U1/aes_core/SB2/n1940 ), 
        .B(\U1/aes_core/SB2/n1939 ), .C(\U1/aes_core/SB2/n1989 ), .D(
        \U1/aes_core/SB2/n1938 ), .Y(\U1/aes_core/SB2/n1941 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1175  ( .A(\U1/aes_core/SB2/n1946 ), .B(
        \U1/aes_core/SB2/n1945 ), .C(\U1/aes_core/SB2/n1944 ), .D(
        \U1/aes_core/SB2/n1943 ), .E(\U1/aes_core/SB2/n1942 ), .F(
        \U1/aes_core/SB2/n1941 ), .Y(\U1/aes_core/SB2/n1987 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1174  ( .A(\U1/aes_core/SB2/n1947 ), .Y(
        \U1/aes_core/SB2/n1951 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1173  ( .A0(\U1/aes_core/SB2/n1949 ), 
        .A1(\U1/aes_core/SB2/n1948 ), .B0(\U1/aes_core/SB2/n1952 ), .B1(
        \U1/aes_core/SB2/n3339 ), .Y(\U1/aes_core/SB2/n1950 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U1172  ( .A0(\U1/aes_core/SB2/n2006 ), 
        .A1(\U1/aes_core/SB2/n3309 ), .B0(\U1/aes_core/SB2/n1951 ), .C0(
        \U1/aes_core/SB2/n1950 ), .Y(\U1/aes_core/SB2/n1961 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1171  ( .A0(\U1/aes_core/SB2/n3276 ), 
        .A1(\U1/aes_core/SB2/n3275 ), .B0(\U1/aes_core/SB2/n3332 ), .Y(
        \U1/aes_core/SB2/n1956 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1170  ( .A0(\U1/aes_core/SB2/n1952 ), 
        .A1(\U1/aes_core/SB2/n3268 ), .B0(\U1/aes_core/SB2/n2060 ), .Y(
        \U1/aes_core/SB2/n1955 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1169  ( .A(\U1/aes_core/SB2/n1956 ), .B(
        \U1/aes_core/SB2/n1955 ), .C(\U1/aes_core/SB2/n1954 ), .D(
        \U1/aes_core/SB2/n1953 ), .Y(\U1/aes_core/SB2/n1960 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1168  ( .A(\U1/aes_core/SB2/n3325 ), .B(
        \U1/aes_core/SB2/n3334 ), .Y(\U1/aes_core/SB2/n1958 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1167  ( .A(\U1/aes_core/SB2/n3331 ), .B(
        \U1/aes_core/SB2/n3333 ), .Y(\U1/aes_core/SB2/n1957 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1166  ( .A(\U1/aes_core/SB2/n1976 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n3310 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1165  ( .A0(\U1/aes_core/SB2/n1958 ), 
        .A1(\U1/aes_core/SB2/n2070 ), .B0(\U1/aes_core/SB2/n1957 ), .B1(
        \U1/aes_core/SB2/n2008 ), .C0(\U1/aes_core/SB2/n3310 ), .C1(
        \U1/aes_core/SB2/n2039 ), .Y(\U1/aes_core/SB2/n1959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1164  ( .A(\U1/aes_core/SB2/n2000 ), .B(
        \U1/aes_core/SB2/n1987 ), .C(\U1/aes_core/SB2/n1962 ), .D(
        \U1/aes_core/SB2/n1961 ), .E(\U1/aes_core/SB2/n1960 ), .F(
        \U1/aes_core/SB2/n1959 ), .Y(\U1/aes_core/sb2 [12]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1163  ( .A(\U1/aes_core/SB2/n3300 ), .B(
        \U1/aes_core/SB2/n3297 ), .Y(\U1/aes_core/SB2/n2025 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U1162  ( .A1N(\U1/aes_core/SB2/n3306 ), 
        .A0(\U1/aes_core/SB2/n3279 ), .B0(\U1/aes_core/SB2/n3344 ), .Y(
        \U1/aes_core/SB2/n1971 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1161  ( .A(\U1/aes_core/SB2/n2053 ), .B(
        \U1/aes_core/SB2/n3268 ), .Y(\U1/aes_core/SB2/n1963 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1160  ( .A0(\U1/aes_core/SB2/n2070 ), 
        .A1(\U1/aes_core/SB2/n3302 ), .B0(\U1/aes_core/SB2/n1963 ), .B1(
        \U1/aes_core/SB2/n3281 ), .C0(\U1/aes_core/SB2/n3297 ), .C1(
        \U1/aes_core/SB2/n3278 ), .Y(\U1/aes_core/SB2/n1970 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1159  ( .A(\U1/aes_core/SB2/n3327 ), .B(
        \U1/aes_core/SB2/n2019 ), .Y(\U1/aes_core/SB2/n2043 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1158  ( .A(\U1/aes_core/SB2/n3299 ), .B(
        \U1/aes_core/SB2/n3282 ), .Y(\U1/aes_core/SB2/n3266 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1157  ( .AN(\U1/aes_core/SB2/n1965 ), 
        .B(\U1/aes_core/SB2/n1964 ), .C(\U1/aes_core/SB2/n2043 ), .D(
        \U1/aes_core/SB2/n3266 ), .Y(\U1/aes_core/SB2/n1969 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1156  ( .A(\U1/aes_core/SB2/n3269 ), .B(
        \U1/aes_core/SB2/n3330 ), .Y(\U1/aes_core/SB2/n3313 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1155  ( .AN(\U1/aes_core/SB2/n1967 ), 
        .B(\U1/aes_core/SB2/n1966 ), .C(\U1/aes_core/SB2/n3313 ), .Y(
        \U1/aes_core/SB2/n1968 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1154  ( .A(\U1/aes_core/SB2/n2025 ), .B(
        \U1/aes_core/SB2/n1972 ), .C(\U1/aes_core/SB2/n1971 ), .D(
        \U1/aes_core/SB2/n1970 ), .E(\U1/aes_core/SB2/n1969 ), .F(
        \U1/aes_core/SB2/n1968 ), .Y(\U1/aes_core/SB2/n2001 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1153  ( .A(\U1/aes_core/SB2/n1973 ), .Y(
        \U1/aes_core/SB2/n1975 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1152  ( .A0(\U1/aes_core/SB2/n3322 ), 
        .A1(\U1/aes_core/SB2/n2058 ), .B0(\U1/aes_core/SB2/n2060 ), .B1(
        \U1/aes_core/SB2/n3327 ), .Y(\U1/aes_core/SB2/n1974 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U1151  ( .A0(\U1/aes_core/SB2/n3344 ), 
        .A1(\U1/aes_core/SB2/n3346 ), .B0(\U1/aes_core/SB2/n1975 ), .C0(
        \U1/aes_core/SB2/n1974 ), .Y(\U1/aes_core/SB2/n1986 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1150  ( .A0(\U1/aes_core/SB2/n3324 ), 
        .A1(\U1/aes_core/SB2/n3322 ), .B0(\U1/aes_core/SB2/n2019 ), .Y(
        \U1/aes_core/SB2/n1979 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1149  ( .A0(\U1/aes_core/SB2/n3325 ), 
        .A1(\U1/aes_core/SB2/n3339 ), .B0(\U1/aes_core/SB2/n1976 ), .Y(
        \U1/aes_core/SB2/n1978 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1148  ( .AN(\U1/aes_core/SB2/n1980 ), 
        .B(\U1/aes_core/SB2/n1979 ), .C(\U1/aes_core/SB2/n1978 ), .D(
        \U1/aes_core/SB2/n1977 ), .Y(\U1/aes_core/SB2/n1985 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1147  ( .A0(\U1/aes_core/SB2/n3332 ), 
        .A1(\U1/aes_core/SB2/n3329 ), .B0(\U1/aes_core/SB2/n3333 ), .Y(
        \U1/aes_core/SB2/n1982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1146  ( .A(\U1/aes_core/SB2/n2017 ), .B(
        \U1/aes_core/SB2/n3302 ), .Y(\U1/aes_core/SB2/n3341 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1145  ( .A0(\U1/aes_core/SB2/n3307 ), 
        .A1(\U1/aes_core/SB2/n3341 ), .B0(\U1/aes_core/SB2/n2054 ), .B1(
        \U1/aes_core/SB2/n3305 ), .Y(\U1/aes_core/SB2/n1981 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U1144  ( .A0(\U1/aes_core/SB2/n1983 ), 
        .A1(\U1/aes_core/SB2/n2039 ), .B0(\U1/aes_core/SB2/n1982 ), .C0(
        \U1/aes_core/SB2/n1981 ), .Y(\U1/aes_core/SB2/n1984 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1143  ( .A(\U1/aes_core/SB2/n2001 ), .B(
        \U1/aes_core/SB2/n1988 ), .C(\U1/aes_core/SB2/n1987 ), .D(
        \U1/aes_core/SB2/n1986 ), .E(\U1/aes_core/SB2/n1985 ), .F(
        \U1/aes_core/SB2/n1984 ), .Y(\U1/aes_core/sb2 [13]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1142  ( .A0(\U1/aes_core/SB2/n3343 ), 
        .A1(\U1/aes_core/SB2/n3296 ), .B0(\U1/aes_core/SB2/n3301 ), .B1(
        \U1/aes_core/SB2/n2070 ), .C0(\U1/aes_core/SB2/n1989 ), .Y(
        \U1/aes_core/SB2/n1998 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1141  ( .A0(\U1/aes_core/SB2/n3275 ), 
        .A1(\U1/aes_core/SB2/n2068 ), .B0(\U1/aes_core/SB2/n3322 ), .Y(
        \U1/aes_core/SB2/n1993 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1140  ( .A0(\U1/aes_core/SB2/n2055 ), 
        .A1(\U1/aes_core/SB2/n3299 ), .B0(\U1/aes_core/SB2/n2060 ), .Y(
        \U1/aes_core/SB2/n1992 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1139  ( .A(\U1/aes_core/SB2/n2010 ), .B(
        \U1/aes_core/SB2/n3346 ), .Y(\U1/aes_core/SB2/n3328 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1138  ( .A0(\U1/aes_core/SB2/n3305 ), 
        .A1(\U1/aes_core/SB2/n3268 ), .B0(\U1/aes_core/SB2/n3328 ), .Y(
        \U1/aes_core/SB2/n1991 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1137  ( .A(\U1/aes_core/SB2/n1993 ), .B(
        \U1/aes_core/SB2/n1992 ), .C(\U1/aes_core/SB2/n1991 ), .D(
        \U1/aes_core/SB2/n1990 ), .Y(\U1/aes_core/SB2/n1997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1136  ( .A(\U1/aes_core/SB2/n3343 ), .B(
        \U1/aes_core/SB2/n3344 ), .Y(\U1/aes_core/SB2/n2066 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1135  ( .A(\U1/aes_core/SB2/n3332 ), .B(
        \U1/aes_core/SB2/n2066 ), .Y(\U1/aes_core/SB2/n1994 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1134  ( .A0(\U1/aes_core/SB2/n2057 ), 
        .A1(\U1/aes_core/SB2/n1995 ), .B0(\U1/aes_core/SB2/n1994 ), .B1(
        \U1/aes_core/SB2/n2010 ), .C0(\U1/aes_core/SB2/n2008 ), .C1(
        \U1/aes_core/SB2/n2039 ), .Y(\U1/aes_core/SB2/n1996 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1133  ( .A(\U1/aes_core/SB2/n2001 ), .B(
        \U1/aes_core/SB2/n2000 ), .C(\U1/aes_core/SB2/n1999 ), .D(
        \U1/aes_core/SB2/n1998 ), .E(\U1/aes_core/SB2/n1997 ), .F(
        \U1/aes_core/SB2/n1996 ), .Y(\U1/aes_core/sb2 [14]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1132  ( .A0(\U1/aes_core/SB2/n2002 ), 
        .A1(\U1/aes_core/SB2/n3302 ), .B0(\U1/aes_core/SB2/n2070 ), .Y(
        \U1/aes_core/SB2/n2014 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U1131  ( .A(\U1/aes_core/SB2/n2005 ), .B(
        \U1/aes_core/SB2/n2004 ), .C(\U1/aes_core/SB2/n2003 ), .Y(
        \U1/aes_core/SB2/n2013 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U1130  ( .A(\U1/aes_core/SB2/n2054 ), .B(
        \U1/aes_core/SB2/n2058 ), .C(\U1/aes_core/SB2/n3282 ), .Y(
        \U1/aes_core/SB2/n2007 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1129  ( .A0(\U1/aes_core/SB2/n2009 ), 
        .A1(\U1/aes_core/SB2/n2008 ), .B0(\U1/aes_core/SB2/n2007 ), .B1(
        \U1/aes_core/SB2/n2065 ), .C0(\U1/aes_core/SB2/n2006 ), .C1(
        \U1/aes_core/SB2/n3280 ), .Y(\U1/aes_core/SB2/n2012 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U1128  ( .A0(\U1/aes_core/SB2/n3343 ), 
        .A1(\U1/aes_core/SB2/n2039 ), .B0(\U1/aes_core/SB2/n3344 ), .B1(
        \U1/aes_core/SB2/n2010 ), .Y(\U1/aes_core/SB2/n2011 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1127  ( .A(\U1/aes_core/SB2/n2016 ), .B(
        \U1/aes_core/SB2/n2015 ), .C(\U1/aes_core/SB2/n2014 ), .D(
        \U1/aes_core/SB2/n2013 ), .E(\U1/aes_core/SB2/n2012 ), .F(
        \U1/aes_core/SB2/n2011 ), .Y(\U1/aes_core/SB2/n3352 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U1126  ( .A0(\U1/aes_core/SB2/n3278 ), 
        .A1(\U1/aes_core/SB2/n3347 ), .B0(\U1/aes_core/SB2/n2017 ), .Y(
        \U1/aes_core/SB2/n2033 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB2/U1125  ( .A0(\U1/aes_core/SB2/n2019 ), 
        .A1(\U1/aes_core/SB2/n3269 ), .B0(\U1/aes_core/SB2/n2018 ), .B1(
        \U1/aes_core/SB2/n3329 ), .Y(\U1/aes_core/SB2/n2032 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1124  ( .A0(\U1/aes_core/SB2/n3281 ), 
        .A1(\U1/aes_core/SB2/n3344 ), .B0(\U1/aes_core/SB2/n2021 ), .B1(
        \U1/aes_core/SB2/n2020 ), .C0(\U1/aes_core/SB2/n2039 ), .C1(
        \U1/aes_core/SB2/n2065 ), .Y(\U1/aes_core/SB2/n2031 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1123  ( .A(\U1/aes_core/SB2/n2025 ), .B(
        \U1/aes_core/SB2/n2024 ), .C(\U1/aes_core/SB2/n2023 ), .D(
        \U1/aes_core/SB2/n2022 ), .Y(\U1/aes_core/SB2/n2030 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1122  ( .AN(\U1/aes_core/SB2/n2028 ), 
        .B(\U1/aes_core/SB2/n2027 ), .C(\U1/aes_core/SB2/n2026 ), .Y(
        \U1/aes_core/SB2/n2029 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1121  ( .A(\U1/aes_core/SB2/n2034 ), .B(
        \U1/aes_core/SB2/n2033 ), .C(\U1/aes_core/SB2/n2032 ), .D(
        \U1/aes_core/SB2/n2031 ), .E(\U1/aes_core/SB2/n2030 ), .F(
        \U1/aes_core/SB2/n2029 ), .Y(\U1/aes_core/SB2/n3294 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1120  ( .A0(\U1/aes_core/SB2/n3307 ), 
        .A1(\U1/aes_core/SB2/n3327 ), .B0(\U1/aes_core/SB2/n2054 ), .Y(
        \U1/aes_core/SB2/n2038 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1119  ( .A(\U1/aes_core/SB2/n2038 ), .B(
        \U1/aes_core/SB2/n2037 ), .C(\U1/aes_core/SB2/n2036 ), .D(
        \U1/aes_core/SB2/n2035 ), .Y(\U1/aes_core/SB2/n2051 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1118  ( .A0(\U1/aes_core/SB2/n3301 ), 
        .A1(\U1/aes_core/SB2/n2070 ), .B0(\U1/aes_core/SB2/n3279 ), .B1(
        \U1/aes_core/SB2/n3280 ), .C0(\U1/aes_core/SB2/n3309 ), .C1(
        \U1/aes_core/SB2/n2039 ), .Y(\U1/aes_core/SB2/n2050 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1117  ( .A(\U1/aes_core/SB2/n2043 ), .B(
        \U1/aes_core/SB2/n2042 ), .C(\U1/aes_core/SB2/n2041 ), .D(
        \U1/aes_core/SB2/n2040 ), .Y(\U1/aes_core/SB2/n2049 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U1116  ( .A(\U1/aes_core/SB2/n2047 ), .B(
        \U1/aes_core/SB2/n2046 ), .C(\U1/aes_core/SB2/n2045 ), .D(
        \U1/aes_core/SB2/n2044 ), .Y(\U1/aes_core/SB2/n2048 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1115  ( .A(\U1/aes_core/SB2/n2051 ), .B(
        \U1/aes_core/SB2/n2050 ), .C(\U1/aes_core/SB2/n2049 ), .D(
        \U1/aes_core/SB2/n2048 ), .Y(\U1/aes_core/SB2/n2052 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1114  ( .A(\U1/aes_core/SB2/n2052 ), .Y(
        \U1/aes_core/SB2/n3285 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1113  ( .A0(\U1/aes_core/SB2/n2055 ), 
        .A1(\U1/aes_core/SB2/n3330 ), .B0(\U1/aes_core/SB2/n2054 ), .B1(
        \U1/aes_core/SB2/n2053 ), .Y(\U1/aes_core/SB2/n2056 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U1112  ( .A0(\U1/aes_core/SB2/n2057 ), 
        .A1(\U1/aes_core/SB2/n3309 ), .B0(\U1/aes_core/SB2/n3285 ), .C0(
        \U1/aes_core/SB2/n2056 ), .Y(\U1/aes_core/SB2/n2073 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U1111  ( .A1N(\U1/aes_core/SB2/n2059 ), 
        .A0(\U1/aes_core/SB2/n2058 ), .B0(\U1/aes_core/SB2/n3332 ), .Y(
        \U1/aes_core/SB2/n2063 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1110  ( .A0(\U1/aes_core/SB2/n3327 ), 
        .A1(\U1/aes_core/SB2/n3322 ), .B0(\U1/aes_core/SB2/n2060 ), .Y(
        \U1/aes_core/SB2/n2062 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1109  ( .AN(\U1/aes_core/SB2/n2064 ), 
        .B(\U1/aes_core/SB2/n2063 ), .C(\U1/aes_core/SB2/n2062 ), .D(
        \U1/aes_core/SB2/n2061 ), .Y(\U1/aes_core/SB2/n2072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1108  ( .A(\U1/aes_core/SB2/n2065 ), .B(
        \U1/aes_core/SB2/n3343 ), .Y(\U1/aes_core/SB2/n2067 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1107  ( .A0(\U1/aes_core/SB2/n2068 ), 
        .A1(\U1/aes_core/SB2/n2067 ), .B0(\U1/aes_core/SB2/n3282 ), .B1(
        \U1/aes_core/SB2/n2066 ), .Y(\U1/aes_core/SB2/n2069 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1106  ( .A0(\U1/aes_core/SB2/n3281 ), 
        .A1(\U1/aes_core/SB2/n3347 ), .B0(\U1/aes_core/SB2/n2070 ), .B1(
        \U1/aes_core/SB2/n3342 ), .C0(\U1/aes_core/SB2/n2069 ), .Y(
        \U1/aes_core/SB2/n2071 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U1105  ( .A(\U1/aes_core/SB2/n3352 ), .B(
        \U1/aes_core/SB2/n3294 ), .C(\U1/aes_core/SB2/n2074 ), .D(
        \U1/aes_core/SB2/n2073 ), .E(\U1/aes_core/SB2/n2072 ), .F(
        \U1/aes_core/SB2/n2071 ), .Y(\U1/aes_core/sb2 [15]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1104  ( .A(Dout[55]), .B(Dout[54]), .Y(
        \U1/aes_core/SB2/n2093 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1103  ( .A(Dout[53]), .B(Dout[52]), .Y(
        \U1/aes_core/SB2/n2084 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1102  ( .A(\U1/aes_core/SB2/n2093 ), .B(
        \U1/aes_core/SB2/n2084 ), .Y(\U1/aes_core/SB2/n2157 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1101  ( .A(Dout[49]), .Y(
        \U1/aes_core/SB2/n2078 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1100  ( .A(Dout[48]), .Y(
        \U1/aes_core/SB2/n2075 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1099  ( .A(\U1/aes_core/SB2/n2078 ), .B(
        \U1/aes_core/SB2/n2075 ), .Y(\U1/aes_core/SB2/n2085 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1098  ( .A(Dout[51]), .B(Dout[50]), .Y(
        \U1/aes_core/SB2/n2105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1097  ( .A(\U1/aes_core/SB2/n2085 ), .B(
        \U1/aes_core/SB2/n2105 ), .Y(\U1/aes_core/SB2/n2464 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1096  ( .A(\U1/aes_core/SB2/n2157 ), .B(
        \U1/aes_core/SB2/n2464 ), .Y(\U1/aes_core/SB2/n2246 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U1095  ( .A(Dout[50]), .B(Dout[51]), .Y(
        \U1/aes_core/SB2/n2088 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1094  ( .A(\U1/aes_core/SB2/n2088 ), .B(
        \U1/aes_core/SB2/n2085 ), .Y(\U1/aes_core/SB2/n2402 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1093  ( .A(Dout[55]), .Y(
        \U1/aes_core/SB2/n2081 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1092  ( .A(\U1/aes_core/SB2/n2081 ), .B(
        Dout[54]), .Y(\U1/aes_core/SB2/n2111 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1091  ( .A(\U1/aes_core/SB2/n2111 ), .B(
        \U1/aes_core/SB2/n2084 ), .Y(\U1/aes_core/SB2/n2156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1090  ( .A(\U1/aes_core/SB2/n2402 ), .B(
        \U1/aes_core/SB2/n2156 ), .Y(\U1/aes_core/SB2/n2368 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1089  ( .A(Dout[51]), .Y(
        \U1/aes_core/SB2/n2076 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U1088  ( .A(Dout[50]), .B(
        \U1/aes_core/SB2/n2076 ), .Y(\U1/aes_core/SB2/n2086 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1087  ( .A(\U1/aes_core/SB2/n2085 ), .B(
        \U1/aes_core/SB2/n2086 ), .Y(\U1/aes_core/SB2/n2308 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1086  ( .A(\U1/aes_core/SB2/n2308 ), .Y(
        \U1/aes_core/SB2/n2498 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1085  ( .A(Dout[52]), .Y(
        \U1/aes_core/SB2/n2077 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1084  ( .A(\U1/aes_core/SB2/n2077 ), .B(
        Dout[53]), .Y(\U1/aes_core/SB2/n2092 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1083  ( .A(Dout[54]), .Y(
        \U1/aes_core/SB2/n2080 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1082  ( .A(\U1/aes_core/SB2/n2080 ), .B(
        Dout[55]), .Y(\U1/aes_core/SB2/n2102 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1081  ( .A(\U1/aes_core/SB2/n2092 ), .B(
        \U1/aes_core/SB2/n2102 ), .Y(\U1/aes_core/SB2/n2354 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1080  ( .A(\U1/aes_core/SB2/n2354 ), .Y(
        \U1/aes_core/SB2/n2452 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1079  ( .A(\U1/aes_core/SB2/n2498 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2286 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1078  ( .A(\U1/aes_core/SB2/n2157 ), .Y(
        \U1/aes_core/SB2/n2467 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1077  ( .A(Dout[49]), .B(Dout[48]), .Y(
        \U1/aes_core/SB2/n2089 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1076  ( .A(\U1/aes_core/SB2/n2089 ), .B(
        \U1/aes_core/SB2/n2105 ), .Y(\U1/aes_core/SB2/n2420 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1075  ( .A(\U1/aes_core/SB2/n2420 ), .Y(
        \U1/aes_core/SB2/n2508 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1074  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2508 ), .Y(\U1/aes_core/SB2/n2425 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1073  ( .A(\U1/aes_core/SB2/n2075 ), .B(
        Dout[49]), .Y(\U1/aes_core/SB2/n2104 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1072  ( .A(\U1/aes_core/SB2/n2086 ), .B(
        \U1/aes_core/SB2/n2104 ), .Y(\U1/aes_core/SB2/n2295 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1071  ( .A(\U1/aes_core/SB2/n2295 ), .Y(
        \U1/aes_core/SB2/n2409 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1070  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2264 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U1069  ( .A(\U1/aes_core/SB2/n2286 ), .B(
        \U1/aes_core/SB2/n2425 ), .C(\U1/aes_core/SB2/n2264 ), .Y(
        \U1/aes_core/SB2/n2124 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1068  ( .A(\U1/aes_core/SB2/n2084 ), .B(
        \U1/aes_core/SB2/n2102 ), .Y(\U1/aes_core/SB2/n2353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1067  ( .A(\U1/aes_core/SB2/n2076 ), .B(
        Dout[50]), .Y(\U1/aes_core/SB2/n2095 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1066  ( .A(\U1/aes_core/SB2/n2095 ), .B(
        \U1/aes_core/SB2/n2104 ), .Y(\U1/aes_core/SB2/n2351 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1065  ( .A(\U1/aes_core/SB2/n2353 ), .B(
        \U1/aes_core/SB2/n2351 ), .Y(\U1/aes_core/SB2/n2241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1064  ( .A(\U1/aes_core/SB2/n2156 ), .Y(
        \U1/aes_core/SB2/n2469 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1063  ( .A(Dout[53]), .Y(
        \U1/aes_core/SB2/n2079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1062  ( .A(\U1/aes_core/SB2/n2077 ), .B(
        \U1/aes_core/SB2/n2079 ), .Y(\U1/aes_core/SB2/n2103 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1061  ( .A(\U1/aes_core/SB2/n2093 ), .B(
        \U1/aes_core/SB2/n2103 ), .Y(\U1/aes_core/SB2/n2512 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1060  ( .A(\U1/aes_core/SB2/n2512 ), .Y(
        \U1/aes_core/SB2/n2443 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1059  ( .A(\U1/aes_core/SB2/n2078 ), .B(
        Dout[48]), .Y(\U1/aes_core/SB2/n2094 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1058  ( .A(\U1/aes_core/SB2/n2094 ), .B(
        \U1/aes_core/SB2/n2105 ), .Y(\U1/aes_core/SB2/n2477 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1057  ( .A(\U1/aes_core/SB2/n2477 ), .Y(
        \U1/aes_core/SB2/n2300 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1056  ( .A0(\U1/aes_core/SB2/n2469 ), 
        .A1(\U1/aes_core/SB2/n2443 ), .B0(\U1/aes_core/SB2/n2300 ), .Y(
        \U1/aes_core/SB2/n2083 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1055  ( .A(\U1/aes_core/SB2/n2089 ), .B(
        \U1/aes_core/SB2/n2086 ), .Y(\U1/aes_core/SB2/n2465 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1054  ( .A(\U1/aes_core/SB2/n2465 ), .Y(
        \U1/aes_core/SB2/n2451 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1053  ( .A(\U1/aes_core/SB2/n2079 ), .B(
        Dout[52]), .Y(\U1/aes_core/SB2/n2110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1052  ( .A(\U1/aes_core/SB2/n2102 ), .B(
        \U1/aes_core/SB2/n2110 ), .Y(\U1/aes_core/SB2/n2505 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1051  ( .A(\U1/aes_core/SB2/n2353 ), .B(
        \U1/aes_core/SB2/n2505 ), .Y(\U1/aes_core/SB2/n2219 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1050  ( .A(\U1/aes_core/SB2/n2081 ), .B(
        \U1/aes_core/SB2/n2080 ), .Y(\U1/aes_core/SB2/n2101 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1049  ( .A(\U1/aes_core/SB2/n2092 ), .B(
        \U1/aes_core/SB2/n2101 ), .Y(\U1/aes_core/SB2/n2480 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1048  ( .A(\U1/aes_core/SB2/n2480 ), .Y(
        \U1/aes_core/SB2/n2200 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1047  ( .A0(\U1/aes_core/SB2/n2451 ), 
        .A1(\U1/aes_core/SB2/n2219 ), .B0(\U1/aes_core/SB2/n2200 ), .B1(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2082 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U1046  ( .AN(\U1/aes_core/SB2/n2241 ), 
        .B(\U1/aes_core/SB2/n2083 ), .C(\U1/aes_core/SB2/n2082 ), .Y(
        \U1/aes_core/SB2/n2123 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1045  ( .A(\U1/aes_core/SB2/n2084 ), .B(
        \U1/aes_core/SB2/n2101 ), .Y(\U1/aes_core/SB2/n2370 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1044  ( .A(\U1/aes_core/SB2/n2088 ), .B(
        \U1/aes_core/SB2/n2089 ), .Y(\U1/aes_core/SB2/n2515 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1043  ( .A(\U1/aes_core/SB2/n2111 ), .B(
        \U1/aes_core/SB2/n2092 ), .Y(\U1/aes_core/SB2/n2421 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1042  ( .A(\U1/aes_core/SB2/n2088 ), .B(
        \U1/aes_core/SB2/n2094 ), .Y(\U1/aes_core/SB2/n2418 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1041  ( .A(\U1/aes_core/SB2/n2085 ), .B(
        \U1/aes_core/SB2/n2095 ), .Y(\U1/aes_core/SB2/n2423 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1040  ( .A(\U1/aes_core/SB2/n2423 ), .Y(
        \U1/aes_core/SB2/n2403 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1039  ( .A(\U1/aes_core/SB2/n2505 ), .Y(
        \U1/aes_core/SB2/n2214 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1038  ( .A(\U1/aes_core/SB2/n2086 ), .B(
        \U1/aes_core/SB2/n2094 ), .Y(\U1/aes_core/SB2/n2441 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1037  ( .A(\U1/aes_core/SB2/n2441 ), .Y(
        \U1/aes_core/SB2/n2466 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U1036  ( .A0(\U1/aes_core/SB2/n2403 ), 
        .A1(\U1/aes_core/SB2/n2467 ), .B0(\U1/aes_core/SB2/n2214 ), .B1(
        \U1/aes_core/SB2/n2466 ), .Y(\U1/aes_core/SB2/n2087 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U1035  ( .A0(\U1/aes_core/SB2/n2370 ), 
        .A1(\U1/aes_core/SB2/n2515 ), .B0(\U1/aes_core/SB2/n2421 ), .B1(
        \U1/aes_core/SB2/n2418 ), .C0(\U1/aes_core/SB2/n2087 ), .Y(
        \U1/aes_core/SB2/n2122 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1034  ( .A(\U1/aes_core/SB2/n2423 ), .B(
        \U1/aes_core/SB2/n2370 ), .Y(\U1/aes_core/SB2/n2207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1033  ( .A(\U1/aes_core/SB2/n2418 ), .B(
        \U1/aes_core/SB2/n2353 ), .Y(\U1/aes_core/SB2/n2217 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1032  ( .A(\U1/aes_core/SB2/n2217 ), .Y(
        \U1/aes_core/SB2/n2091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1031  ( .A(\U1/aes_core/SB2/n2088 ), .B(
        \U1/aes_core/SB2/n2104 ), .Y(\U1/aes_core/SB2/n2493 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1030  ( .A(\U1/aes_core/SB2/n2493 ), .Y(
        \U1/aes_core/SB2/n2442 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1029  ( .A(\U1/aes_core/SB2/n2089 ), .B(
        \U1/aes_core/SB2/n2095 ), .Y(\U1/aes_core/SB2/n2478 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1028  ( .A(\U1/aes_core/SB2/n2478 ), .Y(
        \U1/aes_core/SB2/n2489 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U1027  ( .A0(\U1/aes_core/SB2/n2442 ), 
        .A1(\U1/aes_core/SB2/n2489 ), .B0(\U1/aes_core/SB2/n2443 ), .Y(
        \U1/aes_core/SB2/n2090 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1026  ( .A(\U1/aes_core/SB2/n2093 ), .B(
        \U1/aes_core/SB2/n2110 ), .Y(\U1/aes_core/SB2/n2494 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1025  ( .A(\U1/aes_core/SB2/n2494 ), .Y(
        \U1/aes_core/SB2/n2444 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1024  ( .A(\U1/aes_core/SB2/n2444 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2234 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1023  ( .AN(\U1/aes_core/SB2/n2207 ), 
        .B(\U1/aes_core/SB2/n2091 ), .C(\U1/aes_core/SB2/n2090 ), .D(
        \U1/aes_core/SB2/n2234 ), .Y(\U1/aes_core/SB2/n2100 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1022  ( .A(\U1/aes_core/SB2/n2103 ), .B(
        \U1/aes_core/SB2/n2101 ), .Y(\U1/aes_core/SB2/n2514 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1021  ( .A(\U1/aes_core/SB2/n2093 ), .B(
        \U1/aes_core/SB2/n2092 ), .Y(\U1/aes_core/SB2/n2506 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U1020  ( .A0(\U1/aes_core/SB2/n2156 ), 
        .A1(\U1/aes_core/SB2/n2308 ), .B0(\U1/aes_core/SB2/n2514 ), .B1(
        \U1/aes_core/SB2/n2423 ), .C0(\U1/aes_core/SB2/n2506 ), .C1(
        \U1/aes_core/SB2/n2441 ), .Y(\U1/aes_core/SB2/n2099 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1019  ( .A(\U1/aes_core/SB2/n2465 ), .B(
        \U1/aes_core/SB2/n2156 ), .Y(\U1/aes_core/SB2/n2292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1018  ( .A(\U1/aes_core/SB2/n2214 ), .B(
        \U1/aes_core/SB2/n2403 ), .Y(\U1/aes_core/SB2/n2245 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1017  ( .A(\U1/aes_core/SB2/n2466 ), .B(
        \U1/aes_core/SB2/n2467 ), .Y(\U1/aes_core/SB2/n2265 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1016  ( .A(\U1/aes_core/SB2/n2421 ), .Y(
        \U1/aes_core/SB2/n2495 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1015  ( .A(\U1/aes_core/SB2/n2495 ), .B(
        \U1/aes_core/SB2/n2300 ), .Y(\U1/aes_core/SB2/n2303 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1014  ( .AN(\U1/aes_core/SB2/n2292 ), 
        .B(\U1/aes_core/SB2/n2245 ), .C(\U1/aes_core/SB2/n2265 ), .D(
        \U1/aes_core/SB2/n2303 ), .Y(\U1/aes_core/SB2/n2098 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1013  ( .A(\U1/aes_core/SB2/n2111 ), .B(
        \U1/aes_core/SB2/n2103 ), .Y(\U1/aes_core/SB2/n2215 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1012  ( .A(\U1/aes_core/SB2/n2215 ), .B(
        \U1/aes_core/SB2/n2477 ), .Y(\U1/aes_core/SB2/n2394 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1011  ( .A(\U1/aes_core/SB2/n2095 ), .B(
        \U1/aes_core/SB2/n2094 ), .Y(\U1/aes_core/SB2/n2513 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1010  ( .A(\U1/aes_core/SB2/n2480 ), .B(
        \U1/aes_core/SB2/n2513 ), .Y(\U1/aes_core/SB2/n2359 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1009  ( .A(\U1/aes_core/SB2/n2359 ), .Y(
        \U1/aes_core/SB2/n2096 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1008  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2300 ), .Y(\U1/aes_core/SB2/n2378 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1007  ( .A(\U1/aes_core/SB2/n2513 ), .Y(
        \U1/aes_core/SB2/n2496 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1006  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2496 ), .Y(\U1/aes_core/SB2/n2429 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U1005  ( .AN(\U1/aes_core/SB2/n2394 ), 
        .B(\U1/aes_core/SB2/n2096 ), .C(\U1/aes_core/SB2/n2378 ), .D(
        \U1/aes_core/SB2/n2429 ), .Y(\U1/aes_core/SB2/n2097 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U1004  ( .A(\U1/aes_core/SB2/n2100 ), .B(
        \U1/aes_core/SB2/n2099 ), .C(\U1/aes_core/SB2/n2098 ), .D(
        \U1/aes_core/SB2/n2097 ), .Y(\U1/aes_core/SB2/n2196 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1003  ( .A(\U1/aes_core/SB2/n2420 ), .B(
        \U1/aes_core/SB2/n2215 ), .Y(\U1/aes_core/SB2/n2428 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U1002  ( .A(\U1/aes_core/SB2/n2110 ), .B(
        \U1/aes_core/SB2/n2101 ), .Y(\U1/aes_core/SB2/n2311 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U1001  ( .A(\U1/aes_core/SB2/n2402 ), .B(
        \U1/aes_core/SB2/n2311 ), .Y(\U1/aes_core/SB2/n2282 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U1000  ( .A(\U1/aes_core/SB2/n2514 ), .Y(
        \U1/aes_core/SB2/n2470 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U999  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2451 ), .Y(\U1/aes_core/SB2/n2231 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U998  ( .A0(\U1/aes_core/SB2/n2311 ), 
        .A1(\U1/aes_core/SB2/n2513 ), .B0(\U1/aes_core/SB2/n2231 ), .Y(
        \U1/aes_core/SB2/n2109 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U997  ( .A(\U1/aes_core/SB2/n2351 ), .Y(
        \U1/aes_core/SB2/n2446 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U996  ( .A(\U1/aes_core/SB2/n2446 ), .B(
        \U1/aes_core/SB2/n2469 ), .Y(\U1/aes_core/SB2/n2447 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U995  ( .A(\U1/aes_core/SB2/n2469 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2406 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U994  ( .A(\U1/aes_core/SB2/n2103 ), .B(
        \U1/aes_core/SB2/n2102 ), .Y(\U1/aes_core/SB2/n2476 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U993  ( .A(\U1/aes_core/SB2/n2476 ), .Y(
        \U1/aes_core/SB2/n2226 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U992  ( .A(\U1/aes_core/SB2/n2442 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2250 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U991  ( .A(\U1/aes_core/SB2/n2464 ), .Y(
        \U1/aes_core/SB2/n2445 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U990  ( .A(\U1/aes_core/SB2/n2445 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2314 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U989  ( .A(\U1/aes_core/SB2/n2447 ), .B(
        \U1/aes_core/SB2/n2406 ), .C(\U1/aes_core/SB2/n2250 ), .D(
        \U1/aes_core/SB2/n2314 ), .Y(\U1/aes_core/SB2/n2108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U988  ( .A(\U1/aes_core/SB2/n2466 ), .B(
        \U1/aes_core/SB2/n2444 ), .Y(\U1/aes_core/SB2/n2373 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U987  ( .A(\U1/aes_core/SB2/n2508 ), .B(
        \U1/aes_core/SB2/n2444 ), .Y(\U1/aes_core/SB2/n2364 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U986  ( .A(\U1/aes_core/SB2/n2506 ), .Y(
        \U1/aes_core/SB2/n2499 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U985  ( .A(\U1/aes_core/SB2/n2403 ), .B(
        \U1/aes_core/SB2/n2499 ), .Y(\U1/aes_core/SB2/n2211 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U984  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2442 ), .Y(\U1/aes_core/SB2/n2347 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U983  ( .A(\U1/aes_core/SB2/n2373 ), .B(
        \U1/aes_core/SB2/n2364 ), .C(\U1/aes_core/SB2/n2211 ), .D(
        \U1/aes_core/SB2/n2347 ), .Y(\U1/aes_core/SB2/n2107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U982  ( .A(\U1/aes_core/SB2/n2418 ), .Y(
        \U1/aes_core/SB2/n2387 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U981  ( .A(\U1/aes_core/SB2/n2214 ), .B(
        \U1/aes_core/SB2/n2387 ), .Y(\U1/aes_core/SB2/n2198 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U980  ( .A(\U1/aes_core/SB2/n2105 ), .B(
        \U1/aes_core/SB2/n2104 ), .Y(\U1/aes_core/SB2/n2453 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U979  ( .A(\U1/aes_core/SB2/n2453 ), .Y(
        \U1/aes_core/SB2/n2487 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U978  ( .A(\U1/aes_core/SB2/n2214 ), .B(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2262 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U977  ( .A(\U1/aes_core/SB2/n2402 ), .Y(
        \U1/aes_core/SB2/n2510 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U976  ( .A(\U1/aes_core/SB2/n2510 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2297 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U975  ( .A(\U1/aes_core/SB2/n2443 ), .B(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2471 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U974  ( .A(\U1/aes_core/SB2/n2198 ), .B(
        \U1/aes_core/SB2/n2262 ), .C(\U1/aes_core/SB2/n2297 ), .D(
        \U1/aes_core/SB2/n2471 ), .Y(\U1/aes_core/SB2/n2106 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U973  ( .A(\U1/aes_core/SB2/n2428 ), .B(
        \U1/aes_core/SB2/n2282 ), .C(\U1/aes_core/SB2/n2109 ), .D(
        \U1/aes_core/SB2/n2108 ), .E(\U1/aes_core/SB2/n2107 ), .F(
        \U1/aes_core/SB2/n2106 ), .Y(\U1/aes_core/SB2/n2185 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U972  ( .A(\U1/aes_core/SB2/n2185 ), .Y(
        \U1/aes_core/SB2/n2120 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U971  ( .A(\U1/aes_core/SB2/n2478 ), .B(
        \U1/aes_core/SB2/n2311 ), .Y(\U1/aes_core/SB2/n2208 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U970  ( .A(\U1/aes_core/SB2/n2111 ), .B(
        \U1/aes_core/SB2/n2110 ), .Y(\U1/aes_core/SB2/n2475 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U969  ( .A(\U1/aes_core/SB2/n2475 ), .B(
        \U1/aes_core/SB2/n2351 ), .Y(\U1/aes_core/SB2/n2360 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U968  ( .A(\U1/aes_core/SB2/n2360 ), .Y(
        \U1/aes_core/SB2/n2113 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U967  ( .A(\U1/aes_core/SB2/n2353 ), .Y(
        \U1/aes_core/SB2/n2500 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U966  ( .A0(\U1/aes_core/SB2/n2226 ), 
        .A1(\U1/aes_core/SB2/n2500 ), .B0(\U1/aes_core/SB2/n2487 ), .Y(
        \U1/aes_core/SB2/n2112 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U965  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2387 ), .Y(\U1/aes_core/SB2/n2233 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U964  ( .AN(\U1/aes_core/SB2/n2208 ), 
        .B(\U1/aes_core/SB2/n2113 ), .C(\U1/aes_core/SB2/n2112 ), .D(
        \U1/aes_core/SB2/n2233 ), .Y(\U1/aes_core/SB2/n2117 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U963  ( .A0(\U1/aes_core/SB2/n2464 ), 
        .A1(\U1/aes_core/SB2/n2512 ), .B0(\U1/aes_core/SB2/n2370 ), .B1(
        \U1/aes_core/SB2/n2418 ), .C0(\U1/aes_core/SB2/n2477 ), .C1(
        \U1/aes_core/SB2/n2494 ), .Y(\U1/aes_core/SB2/n2116 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U962  ( .A(\U1/aes_core/SB2/n2512 ), .B(
        \U1/aes_core/SB2/n2515 ), .Y(\U1/aes_core/SB2/n2273 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U961  ( .A(\U1/aes_core/SB2/n2500 ), .B(
        \U1/aes_core/SB2/n2442 ), .Y(\U1/aes_core/SB2/n2431 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U960  ( .A(\U1/aes_core/SB2/n2403 ), .B(
        \U1/aes_core/SB2/n2500 ), .Y(\U1/aes_core/SB2/n2365 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U959  ( .A(\U1/aes_core/SB2/n2387 ), .B(
        \U1/aes_core/SB2/n2467 ), .Y(\U1/aes_core/SB2/n2212 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U958  ( .AN(\U1/aes_core/SB2/n2273 ), 
        .B(\U1/aes_core/SB2/n2431 ), .C(\U1/aes_core/SB2/n2365 ), .D(
        \U1/aes_core/SB2/n2212 ), .Y(\U1/aes_core/SB2/n2115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U957  ( .A(\U1/aes_core/SB2/n2510 ), .B(
        \U1/aes_core/SB2/n2495 ), .Y(\U1/aes_core/SB2/n2285 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U956  ( .A(\U1/aes_core/SB2/n2387 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2377 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U955  ( .A(\U1/aes_core/SB2/n2214 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U954  ( .A(\U1/aes_core/SB2/n2446 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2298 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U953  ( .A(\U1/aes_core/SB2/n2285 ), .B(
        \U1/aes_core/SB2/n2377 ), .C(\U1/aes_core/SB2/n2253 ), .D(
        \U1/aes_core/SB2/n2298 ), .Y(\U1/aes_core/SB2/n2114 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U952  ( .A(\U1/aes_core/SB2/n2117 ), .B(
        \U1/aes_core/SB2/n2116 ), .C(\U1/aes_core/SB2/n2115 ), .D(
        \U1/aes_core/SB2/n2114 ), .Y(\U1/aes_core/SB2/n2118 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U951  ( .A(\U1/aes_core/SB2/n2118 ), .Y(
        \U1/aes_core/SB2/n2492 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U950  ( .A(\U1/aes_core/SB2/n2508 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2119 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U949  ( .AN(\U1/aes_core/SB2/n2196 ), 
        .B(\U1/aes_core/SB2/n2120 ), .C(\U1/aes_core/SB2/n2492 ), .D(
        \U1/aes_core/SB2/n2119 ), .Y(\U1/aes_core/SB2/n2121 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U948  ( .A(\U1/aes_core/SB2/n2246 ), .B(
        \U1/aes_core/SB2/n2368 ), .C(\U1/aes_core/SB2/n2124 ), .D(
        \U1/aes_core/SB2/n2123 ), .E(\U1/aes_core/SB2/n2122 ), .F(
        \U1/aes_core/SB2/n2121 ), .Y(\U1/aes_core/SB2/n2175 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U947  ( .A(\U1/aes_core/SB2/n2493 ), .B(
        \U1/aes_core/SB2/n2156 ), .Y(\U1/aes_core/SB2/n2291 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U946  ( .A(\U1/aes_core/SB2/n2443 ), .B(
        \U1/aes_core/SB2/n2510 ), .Y(\U1/aes_core/SB2/n2367 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U945  ( .A(\U1/aes_core/SB2/n2499 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2244 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U944  ( .A(\U1/aes_core/SB2/n2215 ), .Y(
        \U1/aes_core/SB2/n2488 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U943  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2267 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U942  ( .AN(\U1/aes_core/SB2/n2291 ), 
        .B(\U1/aes_core/SB2/n2367 ), .C(\U1/aes_core/SB2/n2244 ), .D(
        \U1/aes_core/SB2/n2267 ), .Y(\U1/aes_core/SB2/n2131 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U941  ( .A(\U1/aes_core/SB2/n2480 ), .B(
        \U1/aes_core/SB2/n2351 ), .Y(\U1/aes_core/SB2/n2393 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U940  ( .A(\U1/aes_core/SB2/n2403 ), .B(
        \U1/aes_core/SB2/n2469 ), .Y(\U1/aes_core/SB2/n2224 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U939  ( .A0(\U1/aes_core/SB2/n2489 ), 
        .A1(\U1/aes_core/SB2/n2409 ), .B0(\U1/aes_core/SB2/n2214 ), .Y(
        \U1/aes_core/SB2/n2125 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U938  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2316 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U937  ( .AN(\U1/aes_core/SB2/n2393 ), 
        .B(\U1/aes_core/SB2/n2224 ), .C(\U1/aes_core/SB2/n2125 ), .D(
        \U1/aes_core/SB2/n2316 ), .Y(\U1/aes_core/SB2/n2126 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U936  ( .A(\U1/aes_core/SB2/n2126 ), .Y(
        \U1/aes_core/SB2/n2130 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U935  ( .A(\U1/aes_core/SB2/n2370 ), .Y(
        \U1/aes_core/SB2/n2490 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U934  ( .A(\U1/aes_core/SB2/n2515 ), .Y(
        \U1/aes_core/SB2/n2410 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U933  ( .A0(\U1/aes_core/SB2/n2510 ), 
        .A1(\U1/aes_core/SB2/n2444 ), .B0(\U1/aes_core/SB2/n2490 ), .B1(
        \U1/aes_core/SB2/n2300 ), .C0(\U1/aes_core/SB2/n2410 ), .C1(
        \U1/aes_core/SB2/n2488 ), .Y(\U1/aes_core/SB2/n2129 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U932  ( .A0(\U1/aes_core/SB2/n2311 ), 
        .A1(\U1/aes_core/SB2/n2493 ), .B0(\U1/aes_core/SB2/n2513 ), .B1(
        \U1/aes_core/SB2/n2514 ), .Y(\U1/aes_core/SB2/n2127 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U931  ( .A0(\U1/aes_core/SB2/n2387 ), 
        .A1(\U1/aes_core/SB2/n2200 ), .B0(\U1/aes_core/SB2/n2443 ), .B1(
        \U1/aes_core/SB2/n2466 ), .C0(\U1/aes_core/SB2/n2127 ), .Y(
        \U1/aes_core/SB2/n2128 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U930  ( .AN(\U1/aes_core/SB2/n2131 ), 
        .B(\U1/aes_core/SB2/n2130 ), .C(\U1/aes_core/SB2/n2129 ), .D(
        \U1/aes_core/SB2/n2128 ), .Y(\U1/aes_core/SB2/n2194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U929  ( .A(\U1/aes_core/SB2/n2514 ), .B(
        \U1/aes_core/SB2/n2351 ), .Y(\U1/aes_core/SB2/n2209 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U928  ( .A0(\U1/aes_core/SB2/n2421 ), 
        .A1(\U1/aes_core/SB2/n2514 ), .B0(\U1/aes_core/SB2/n2453 ), .Y(
        \U1/aes_core/SB2/n2136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U927  ( .A(\U1/aes_core/SB2/n2453 ), .B(
        \U1/aes_core/SB2/n2441 ), .Y(\U1/aes_core/SB2/n2293 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB2/U926  ( .A0(\U1/aes_core/SB2/n2442 ), .A1(
        \U1/aes_core/SB2/n2200 ), .B0(\U1/aes_core/SB2/n2293 ), .B1(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2135 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U925  ( .A0(\U1/aes_core/SB2/n2475 ), 
        .A1(\U1/aes_core/SB2/n2515 ), .B0(\U1/aes_core/SB2/n2215 ), .B1(
        \U1/aes_core/SB2/n2308 ), .C0(\U1/aes_core/SB2/n2477 ), .C1(
        \U1/aes_core/SB2/n2506 ), .Y(\U1/aes_core/SB2/n2134 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U924  ( .A(\U1/aes_core/SB2/n2311 ), .Y(
        \U1/aes_core/SB2/n2404 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U923  ( .A(\U1/aes_core/SB2/n2508 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2430 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U922  ( .A(\U1/aes_core/SB2/n2403 ), .B(
        \U1/aes_core/SB2/n2200 ), .Y(\U1/aes_core/SB2/n2232 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U921  ( .A(\U1/aes_core/SB2/n2214 ), .B(
        \U1/aes_core/SB2/n2446 ), .Y(\U1/aes_core/SB2/n2252 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U920  ( .A(\U1/aes_core/SB2/n2403 ), .B(
        \U1/aes_core/SB2/n2444 ), .Y(\U1/aes_core/SB2/n2376 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U919  ( .A(\U1/aes_core/SB2/n2430 ), .B(
        \U1/aes_core/SB2/n2232 ), .C(\U1/aes_core/SB2/n2252 ), .D(
        \U1/aes_core/SB2/n2376 ), .Y(\U1/aes_core/SB2/n2133 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U918  ( .A(\U1/aes_core/SB2/n2423 ), .B(
        \U1/aes_core/SB2/n2311 ), .Y(\U1/aes_core/SB2/n2274 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U917  ( .A(\U1/aes_core/SB2/n2409 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2284 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U916  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2300 ), .Y(\U1/aes_core/SB2/n2315 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U915  ( .AN(\U1/aes_core/SB2/n2274 ), 
        .B(\U1/aes_core/SB2/n2284 ), .C(\U1/aes_core/SB2/n2315 ), .Y(
        \U1/aes_core/SB2/n2132 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U914  ( .A(\U1/aes_core/SB2/n2209 ), .B(
        \U1/aes_core/SB2/n2136 ), .C(\U1/aes_core/SB2/n2135 ), .D(
        \U1/aes_core/SB2/n2134 ), .E(\U1/aes_core/SB2/n2133 ), .F(
        \U1/aes_core/SB2/n2132 ), .Y(\U1/aes_core/SB2/n2521 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U913  ( .A0(\U1/aes_core/SB2/n2214 ), 
        .A1(\U1/aes_core/SB2/n2467 ), .B0(\U1/aes_core/SB2/n2498 ), .Y(
        \U1/aes_core/SB2/n2137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U912  ( .A(\U1/aes_core/SB2/n2200 ), .B(
        \U1/aes_core/SB2/n2300 ), .Y(\U1/aes_core/SB2/n2362 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U911  ( .A(\U1/aes_core/SB2/n2442 ), .B(
        \U1/aes_core/SB2/n2490 ), .Y(\U1/aes_core/SB2/n2229 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U910  ( .A(\U1/aes_core/SB2/n2490 ), .B(
        \U1/aes_core/SB2/n2446 ), .Y(\U1/aes_core/SB2/n2280 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U909  ( .A(\U1/aes_core/SB2/n2137 ), .B(
        \U1/aes_core/SB2/n2362 ), .C(\U1/aes_core/SB2/n2229 ), .D(
        \U1/aes_core/SB2/n2280 ), .Y(\U1/aes_core/SB2/n2141 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U908  ( .A0(\U1/aes_core/SB2/n2493 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2215 ), .B1(
        \U1/aes_core/SB2/n2465 ), .C0(\U1/aes_core/SB2/n2494 ), .C1(
        \U1/aes_core/SB2/n2351 ), .Y(\U1/aes_core/SB2/n2140 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U907  ( .A(\U1/aes_core/SB2/n2445 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2261 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U906  ( .A(\U1/aes_core/SB2/n2444 ), .B(
        \U1/aes_core/SB2/n2496 ), .Y(\U1/aes_core/SB2/n2426 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U905  ( .A(\U1/aes_core/SB2/n2444 ), .B(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U904  ( .A(\U1/aes_core/SB2/n2499 ), .B(
        \U1/aes_core/SB2/n2489 ), .Y(\U1/aes_core/SB2/n2210 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U903  ( .A(\U1/aes_core/SB2/n2261 ), .B(
        \U1/aes_core/SB2/n2426 ), .C(\U1/aes_core/SB2/n2248 ), .D(
        \U1/aes_core/SB2/n2210 ), .Y(\U1/aes_core/SB2/n2139 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U902  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2348 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U901  ( .A(\U1/aes_core/SB2/n2508 ), .B(
        \U1/aes_core/SB2/n2469 ), .Y(\U1/aes_core/SB2/n2296 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U900  ( .A(\U1/aes_core/SB2/n2498 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2372 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U899  ( .A(\U1/aes_core/SB2/n2226 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2197 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U898  ( .A(\U1/aes_core/SB2/n2348 ), .B(
        \U1/aes_core/SB2/n2296 ), .C(\U1/aes_core/SB2/n2372 ), .D(
        \U1/aes_core/SB2/n2197 ), .Y(\U1/aes_core/SB2/n2138 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U897  ( .A(\U1/aes_core/SB2/n2141 ), .B(
        \U1/aes_core/SB2/n2140 ), .C(\U1/aes_core/SB2/n2139 ), .D(
        \U1/aes_core/SB2/n2138 ), .Y(\U1/aes_core/SB2/n2183 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U896  ( .A(\U1/aes_core/SB2/n2175 ), .B(
        \U1/aes_core/SB2/n2194 ), .C(\U1/aes_core/SB2/n2521 ), .D(
        \U1/aes_core/SB2/n2183 ), .Y(\U1/aes_core/SB2/n2150 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U895  ( .A(\U1/aes_core/SB2/n2475 ), .Y(
        \U1/aes_core/SB2/n2399 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U894  ( .A0(\U1/aes_core/SB2/n2351 ), 
        .A1(\U1/aes_core/SB2/n2157 ), .B0(\U1/aes_core/SB2/n2295 ), .B1(
        \U1/aes_core/SB2/n2506 ), .Y(\U1/aes_core/SB2/n2142 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U893  ( .A0(\U1/aes_core/SB2/n2399 ), 
        .A1(\U1/aes_core/SB2/n2451 ), .B0(\U1/aes_core/SB2/n2500 ), .B1(
        \U1/aes_core/SB2/n2508 ), .C0(\U1/aes_core/SB2/n2142 ), .Y(
        \U1/aes_core/SB2/n2149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U892  ( .A(\U1/aes_core/SB2/n2420 ), .B(
        \U1/aes_core/SB2/n2423 ), .Y(\U1/aes_core/SB2/n2419 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U891  ( .A0(\U1/aes_core/SB2/n2354 ), 
        .A1(\U1/aes_core/SB2/n2423 ), .B0(\U1/aes_core/SB2/n2311 ), .B1(
        \U1/aes_core/SB2/n2464 ), .Y(\U1/aes_core/SB2/n2143 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U890  ( .A0(\U1/aes_core/SB2/n2226 ), 
        .A1(\U1/aes_core/SB2/n2419 ), .B0(\U1/aes_core/SB2/n2470 ), .B1(
        \U1/aes_core/SB2/n2489 ), .C0(\U1/aes_core/SB2/n2143 ), .Y(
        \U1/aes_core/SB2/n2148 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U889  ( .A(\U1/aes_core/SB2/n2494 ), .B(
        \U1/aes_core/SB2/n2353 ), .Y(\U1/aes_core/SB2/n2146 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U888  ( .A(\U1/aes_core/SB2/n2444 ), .B(
        \U1/aes_core/SB2/n2469 ), .Y(\U1/aes_core/SB2/n2411 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U887  ( .A(\U1/aes_core/SB2/n2411 ), .Y(
        \U1/aes_core/SB2/n2145 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U886  ( .A(\U1/aes_core/SB2/n2402 ), .B(
        \U1/aes_core/SB2/n2475 ), .Y(\U1/aes_core/SB2/n2258 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U885  ( .A(\U1/aes_core/SB2/n2480 ), .B(
        \U1/aes_core/SB2/n2478 ), .Y(\U1/aes_core/SB2/n2436 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U883  ( .A(\U1/aes_core/SB2/n2451 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2268 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U881  ( .A0(\U1/aes_core/SB2/n2410 ), 
        .A1(\U1/aes_core/SB2/n2146 ), .B0(\U1/aes_core/SB2/n2387 ), .B1(
        \U1/aes_core/SB2/n2145 ), .C0(\U1/aes_core/SB2/n2144 ), .Y(
        \U1/aes_core/SB2/n2147 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U880  ( .AN(\U1/aes_core/SB2/n2150 ), 
        .B(\U1/aes_core/SB2/n2149 ), .C(\U1/aes_core/SB2/n2148 ), .D(
        \U1/aes_core/SB2/n2147 ), .Y(\U1/aes_core/sb2 [16]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U879  ( .A(\U1/aes_core/SB2/n2423 ), .B(
        \U1/aes_core/SB2/n2215 ), .Y(\U1/aes_core/SB2/n2275 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U878  ( .A(\U1/aes_core/SB2/n2370 ), .B(
        \U1/aes_core/SB2/n2420 ), .Y(\U1/aes_core/SB2/n2235 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U877  ( .A(\U1/aes_core/SB2/n2387 ), .B(
        \U1/aes_core/SB2/n2498 ), .Y(\U1/aes_core/SB2/n2369 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U876  ( .A0(\U1/aes_core/SB2/n2369 ), 
        .A1(\U1/aes_core/SB2/n2423 ), .B0(\U1/aes_core/SB2/n2512 ), .Y(
        \U1/aes_core/SB2/n2155 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U875  ( .A(\U1/aes_core/SB2/n2451 ), .B(
        \U1/aes_core/SB2/n2499 ), .Y(\U1/aes_core/SB2/n2251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U874  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2451 ), .Y(\U1/aes_core/SB2/n2375 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U873  ( .A(\U1/aes_core/SB2/n2496 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2283 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U872  ( .A(\U1/aes_core/SB2/n2251 ), .B(
        \U1/aes_core/SB2/n2375 ), .C(\U1/aes_core/SB2/n2283 ), .Y(
        \U1/aes_core/SB2/n2154 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U871  ( .A(\U1/aes_core/SB2/n2451 ), .B(
        \U1/aes_core/SB2/n2510 ), .Y(\U1/aes_core/SB2/n2310 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U870  ( .A(\U1/aes_core/SB2/n2496 ), .B(
        \U1/aes_core/SB2/n2487 ), .C(\U1/aes_core/SB2/n2508 ), .Y(
        \U1/aes_core/SB2/n2151 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U869  ( .A0(\U1/aes_core/SB2/n2310 ), 
        .A1(\U1/aes_core/SB2/n2476 ), .B0(\U1/aes_core/SB2/n2151 ), .B1(
        \U1/aes_core/SB2/n2506 ), .C0(\U1/aes_core/SB2/n2370 ), .C1(
        \U1/aes_core/SB2/n2402 ), .Y(\U1/aes_core/SB2/n2153 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U868  ( .A0(\U1/aes_core/SB2/n2477 ), 
        .A1(\U1/aes_core/SB2/n2505 ), .B0(\U1/aes_core/SB2/n2478 ), .B1(
        \U1/aes_core/SB2/n2475 ), .Y(\U1/aes_core/SB2/n2152 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U867  ( .A(\U1/aes_core/SB2/n2275 ), .B(
        \U1/aes_core/SB2/n2235 ), .C(\U1/aes_core/SB2/n2155 ), .D(
        \U1/aes_core/SB2/n2154 ), .E(\U1/aes_core/SB2/n2153 ), .F(
        \U1/aes_core/SB2/n2152 ), .Y(\U1/aes_core/SB2/n2520 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U866  ( .A(\U1/aes_core/SB2/n2351 ), .B(
        \U1/aes_core/SB2/n2311 ), .Y(\U1/aes_core/SB2/n2201 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U865  ( .A0(\U1/aes_core/SB2/n2351 ), 
        .A1(\U1/aes_core/SB2/n2441 ), .B0(\U1/aes_core/SB2/n2215 ), .Y(
        \U1/aes_core/SB2/n2162 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U864  ( .A(\U1/aes_core/SB2/n2445 ), .B(
        \U1/aes_core/SB2/n2451 ), .Y(\U1/aes_core/SB2/n2203 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U863  ( .A0(\U1/aes_core/SB2/n2308 ), 
        .A1(\U1/aes_core/SB2/n2480 ), .B0(\U1/aes_core/SB2/n2203 ), .B1(
        \U1/aes_core/SB2/n2494 ), .Y(\U1/aes_core/SB2/n2161 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U862  ( .A0(\U1/aes_core/SB2/n2295 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2464 ), .B1(
        \U1/aes_core/SB2/n2370 ), .C0(\U1/aes_core/SB2/n2478 ), .C1(
        \U1/aes_core/SB2/n2421 ), .Y(\U1/aes_core/SB2/n2160 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U861  ( .A(\U1/aes_core/SB2/n2513 ), .B(
        \U1/aes_core/SB2/n2156 ), .Y(\U1/aes_core/SB2/n2259 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U860  ( .A(\U1/aes_core/SB2/n2500 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2266 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U859  ( .A(\U1/aes_core/SB2/n2442 ), .B(
        \U1/aes_core/SB2/n2495 ), .Y(\U1/aes_core/SB2/n2276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U858  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2510 ), .Y(\U1/aes_core/SB2/n2405 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U857  ( .AN(\U1/aes_core/SB2/n2259 ), 
        .B(\U1/aes_core/SB2/n2266 ), .C(\U1/aes_core/SB2/n2276 ), .D(
        \U1/aes_core/SB2/n2405 ), .Y(\U1/aes_core/SB2/n2159 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U856  ( .A(\U1/aes_core/SB2/n2402 ), .B(
        \U1/aes_core/SB2/n2157 ), .Y(\U1/aes_core/SB2/n2384 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U855  ( .A(\U1/aes_core/SB2/n2480 ), .B(
        \U1/aes_core/SB2/n2464 ), .Y(\U1/aes_core/SB2/n2437 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U853  ( .A(\U1/aes_core/SB2/n2200 ), .B(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2225 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U851  ( .A(\U1/aes_core/SB2/n2201 ), .B(
        \U1/aes_core/SB2/n2162 ), .C(\U1/aes_core/SB2/n2161 ), .D(
        \U1/aes_core/SB2/n2160 ), .E(\U1/aes_core/SB2/n2159 ), .F(
        \U1/aes_core/SB2/n2158 ), .Y(\U1/aes_core/SB2/n2195 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U850  ( .A(\U1/aes_core/SB2/n2418 ), .B(
        \U1/aes_core/SB2/n2215 ), .Y(\U1/aes_core/SB2/n2213 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U849  ( .A(\U1/aes_core/SB2/n2370 ), .B(
        \U1/aes_core/SB2/n2295 ), .Y(\U1/aes_core/SB2/n2450 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U848  ( .A(\U1/aes_core/SB2/n2351 ), .B(
        \U1/aes_core/SB2/n2421 ), .Y(\U1/aes_core/SB2/n2263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U847  ( .A(\U1/aes_core/SB2/n2515 ), .B(
        \U1/aes_core/SB2/n2421 ), .Y(\U1/aes_core/SB2/n2278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U846  ( .A(\U1/aes_core/SB2/n2446 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2363 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U845  ( .A(\U1/aes_core/SB2/n2496 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U844  ( .A(\U1/aes_core/SB2/n2500 ), .B(
        \U1/aes_core/SB2/n2496 ), .Y(\U1/aes_core/SB2/n2349 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U843  ( .A(\U1/aes_core/SB2/n2410 ), .B(
        \U1/aes_core/SB2/n2467 ), .Y(\U1/aes_core/SB2/n2249 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U842  ( .A(\U1/aes_core/SB2/n2363 ), .B(
        \U1/aes_core/SB2/n2230 ), .C(\U1/aes_core/SB2/n2349 ), .D(
        \U1/aes_core/SB2/n2249 ), .Y(\U1/aes_core/SB2/n2166 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U841  ( .A(\U1/aes_core/SB2/n2515 ), .B(
        \U1/aes_core/SB2/n2311 ), .Y(\U1/aes_core/SB2/n2299 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U840  ( .A(\U1/aes_core/SB2/n2514 ), .B(
        \U1/aes_core/SB2/n2295 ), .Y(\U1/aes_core/SB2/n2424 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U839  ( .A(\U1/aes_core/SB2/n2441 ), .B(
        \U1/aes_core/SB2/n2480 ), .Y(\U1/aes_core/SB2/n2374 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U838  ( .A(\U1/aes_core/SB2/n2402 ), .B(
        \U1/aes_core/SB2/n2480 ), .Y(\U1/aes_core/SB2/n2199 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U837  ( .A0(\U1/aes_core/SB2/n2480 ), 
        .A1(\U1/aes_core/SB2/n2515 ), .B0(\U1/aes_core/SB2/n2311 ), .B1(
        \U1/aes_core/SB2/n2441 ), .Y(\U1/aes_core/SB2/n2164 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U836  ( .A0(\U1/aes_core/SB2/n2295 ), 
        .A1(\U1/aes_core/SB2/n2512 ), .B0(\U1/aes_core/SB2/n2308 ), .B1(
        \U1/aes_core/SB2/n2370 ), .Y(\U1/aes_core/SB2/n2163 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U835  ( .A(\U1/aes_core/SB2/n2299 ), .B(
        \U1/aes_core/SB2/n2424 ), .C(\U1/aes_core/SB2/n2374 ), .D(
        \U1/aes_core/SB2/n2199 ), .E(\U1/aes_core/SB2/n2164 ), .F(
        \U1/aes_core/SB2/n2163 ), .Y(\U1/aes_core/SB2/n2165 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U834  ( .A(\U1/aes_core/SB2/n2213 ), .B(
        \U1/aes_core/SB2/n2450 ), .C(\U1/aes_core/SB2/n2263 ), .D(
        \U1/aes_core/SB2/n2278 ), .E(\U1/aes_core/SB2/n2166 ), .F(
        \U1/aes_core/SB2/n2165 ), .Y(\U1/aes_core/SB2/n2184 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U833  ( .A0(\U1/aes_core/SB2/n2446 ), 
        .A1(\U1/aes_core/SB2/n2443 ), .B0(\U1/aes_core/SB2/n2499 ), .B1(
        \U1/aes_core/SB2/n2387 ), .C0(\U1/aes_core/SB2/n2184 ), .Y(
        \U1/aes_core/SB2/n2167 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U832  ( .A(\U1/aes_core/SB2/n2167 ), .Y(
        \U1/aes_core/SB2/n2174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U831  ( .A(\U1/aes_core/SB2/n2478 ), .B(
        \U1/aes_core/SB2/n2441 ), .Y(\U1/aes_core/SB2/n2468 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U830  ( .A0(\U1/aes_core/SB2/n2445 ), 
        .A1(\U1/aes_core/SB2/n2468 ), .B0(\U1/aes_core/SB2/n2500 ), .Y(
        \U1/aes_core/SB2/n2170 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U829  ( .A0(\U1/aes_core/SB2/n2410 ), 
        .A1(\U1/aes_core/SB2/n2489 ), .B0(\U1/aes_core/SB2/n2452 ), .Y(
        \U1/aes_core/SB2/n2169 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U828  ( .A0(\U1/aes_core/SB2/n2409 ), 
        .A1(\U1/aes_core/SB2/n2451 ), .B0(\U1/aes_core/SB2/n2495 ), .Y(
        \U1/aes_core/SB2/n2168 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U827  ( .A(\U1/aes_core/SB2/n2442 ), .B(
        \U1/aes_core/SB2/n2488 ), .Y(\U1/aes_core/SB2/n2242 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U826  ( .A(\U1/aes_core/SB2/n2170 ), .B(
        \U1/aes_core/SB2/n2169 ), .C(\U1/aes_core/SB2/n2168 ), .D(
        \U1/aes_core/SB2/n2242 ), .Y(\U1/aes_core/SB2/n2173 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U825  ( .A(\U1/aes_core/SB2/n2487 ), .B(
        \U1/aes_core/SB2/n2403 ), .Y(\U1/aes_core/SB2/n2457 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB2/U824  ( .A(\U1/aes_core/SB2/n2457 ), .B(
        \U1/aes_core/SB2/n2477 ), .C(\U1/aes_core/SB2/n2464 ), .Y(
        \U1/aes_core/SB2/n2171 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U823  ( .A0(\U1/aes_core/SB2/n2441 ), 
        .A1(\U1/aes_core/SB2/n2514 ), .B0(\U1/aes_core/SB2/n2171 ), .B1(
        \U1/aes_core/SB2/n2475 ), .C0(\U1/aes_core/SB2/n2513 ), .C1(
        \U1/aes_core/SB2/n2505 ), .Y(\U1/aes_core/SB2/n2172 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U822  ( .A(\U1/aes_core/SB2/n2520 ), .B(
        \U1/aes_core/SB2/n2195 ), .C(\U1/aes_core/SB2/n2175 ), .D(
        \U1/aes_core/SB2/n2174 ), .E(\U1/aes_core/SB2/n2173 ), .F(
        \U1/aes_core/SB2/n2172 ), .Y(\U1/aes_core/sb2 [17]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U821  ( .A0(\U1/aes_core/SB2/n2469 ), 
        .A1(\U1/aes_core/SB2/n2489 ), .B0(\U1/aes_core/SB2/n2510 ), .B1(
        \U1/aes_core/SB2/n2500 ), .Y(\U1/aes_core/SB2/n2176 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U820  ( .A0(\U1/aes_core/SB2/n2420 ), 
        .A1(\U1/aes_core/SB2/n2514 ), .B0(\U1/aes_core/SB2/n2370 ), .B1(
        \U1/aes_core/SB2/n2441 ), .C0(\U1/aes_core/SB2/n2176 ), .Y(
        \U1/aes_core/SB2/n2182 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U819  ( .A(\U1/aes_core/SB2/n2495 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2279 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U818  ( .A(\U1/aes_core/SB2/n2469 ), .B(
        \U1/aes_core/SB2/n2445 ), .Y(\U1/aes_core/SB2/n2260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U817  ( .A(\U1/aes_core/SB2/n2489 ), .B(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2228 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U816  ( .A(\U1/aes_core/SB2/n2409 ), .B(
        \U1/aes_core/SB2/n2452 ), .Y(\U1/aes_core/SB2/n2247 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U815  ( .A(\U1/aes_core/SB2/n2279 ), .B(
        \U1/aes_core/SB2/n2260 ), .C(\U1/aes_core/SB2/n2228 ), .D(
        \U1/aes_core/SB2/n2247 ), .Y(\U1/aes_core/SB2/n2181 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U814  ( .A(\U1/aes_core/SB2/n2515 ), .B(
        \U1/aes_core/SB2/n2493 ), .Y(\U1/aes_core/SB2/n2398 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U813  ( .A0(\U1/aes_core/SB2/n2446 ), 
        .A1(\U1/aes_core/SB2/n2398 ), .B0(\U1/aes_core/SB2/n2499 ), .Y(
        \U1/aes_core/SB2/n2179 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U812  ( .A0(\U1/aes_core/SB2/n2496 ), 
        .A1(\U1/aes_core/SB2/n2387 ), .B0(\U1/aes_core/SB2/n2399 ), .Y(
        \U1/aes_core/SB2/n2178 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U811  ( .A0(\U1/aes_core/SB2/n2404 ), 
        .A1(\U1/aes_core/SB2/n2444 ), .B0(\U1/aes_core/SB2/n2498 ), .Y(
        \U1/aes_core/SB2/n2177 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U810  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2496 ), .Y(\U1/aes_core/SB2/n2371 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U809  ( .A(\U1/aes_core/SB2/n2179 ), .B(
        \U1/aes_core/SB2/n2178 ), .C(\U1/aes_core/SB2/n2177 ), .D(
        \U1/aes_core/SB2/n2371 ), .Y(\U1/aes_core/SB2/n2180 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U808  ( .A(\U1/aes_core/SB2/n2185 ), .B(
        \U1/aes_core/SB2/n2184 ), .C(\U1/aes_core/SB2/n2183 ), .D(
        \U1/aes_core/SB2/n2182 ), .E(\U1/aes_core/SB2/n2181 ), .F(
        \U1/aes_core/SB2/n2180 ), .Y(\U1/aes_core/SB2/n2519 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U807  ( .A0(\U1/aes_core/SB2/n2300 ), 
        .A1(\U1/aes_core/SB2/n2500 ), .B0(\U1/aes_core/SB2/n2508 ), .B1(
        \U1/aes_core/SB2/n2443 ), .C0(\U1/aes_core/SB2/n2519 ), .Y(
        \U1/aes_core/SB2/n2186 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U806  ( .A(\U1/aes_core/SB2/n2186 ), .Y(
        \U1/aes_core/SB2/n2193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U805  ( .A(\U1/aes_core/SB2/n2452 ), .B(
        \U1/aes_core/SB2/n2214 ), .Y(\U1/aes_core/SB2/n2361 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U804  ( .A1N(\U1/aes_core/SB2/n2361 ), 
        .A0(\U1/aes_core/SB2/n2470 ), .B0(\U1/aes_core/SB2/n2442 ), .Y(
        \U1/aes_core/SB2/n2189 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U803  ( .A0(\U1/aes_core/SB2/n2410 ), 
        .A1(\U1/aes_core/SB2/n2293 ), .B0(\U1/aes_core/SB2/n2469 ), .Y(
        \U1/aes_core/SB2/n2188 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U802  ( .A0(\U1/aes_core/SB2/n2496 ), 
        .A1(\U1/aes_core/SB2/n2451 ), .B0(\U1/aes_core/SB2/n2490 ), .Y(
        \U1/aes_core/SB2/n2187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U801  ( .A(\U1/aes_core/SB2/n2467 ), .B(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2243 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U800  ( .A(\U1/aes_core/SB2/n2189 ), .B(
        \U1/aes_core/SB2/n2188 ), .C(\U1/aes_core/SB2/n2187 ), .D(
        \U1/aes_core/SB2/n2243 ), .Y(\U1/aes_core/SB2/n2192 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U799  ( .A(\U1/aes_core/SB2/n2466 ), .B(
        \U1/aes_core/SB2/n2498 ), .Y(\U1/aes_core/SB2/n2497 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U798  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2444 ), .Y(\U1/aes_core/SB2/n2190 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U797  ( .A0(\U1/aes_core/SB2/n2497 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2190 ), .B1(
        \U1/aes_core/SB2/n2478 ), .C0(\U1/aes_core/SB2/n2421 ), .C1(
        \U1/aes_core/SB2/n2423 ), .Y(\U1/aes_core/SB2/n2191 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U796  ( .A(\U1/aes_core/SB2/n2196 ), .B(
        \U1/aes_core/SB2/n2195 ), .C(\U1/aes_core/SB2/n2194 ), .D(
        \U1/aes_core/SB2/n2193 ), .E(\U1/aes_core/SB2/n2192 ), .F(
        \U1/aes_core/SB2/n2191 ), .Y(\U1/aes_core/sb2 [18]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U795  ( .A(\U1/aes_core/SB2/n2300 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2502 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U794  ( .AN(\U1/aes_core/SB2/n2199 ), 
        .B(\U1/aes_core/SB2/n2198 ), .C(\U1/aes_core/SB2/n2197 ), .D(
        \U1/aes_core/SB2/n2502 ), .Y(\U1/aes_core/SB2/n2206 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U793  ( .A0(\U1/aes_core/SB2/n2200 ), 
        .A1(\U1/aes_core/SB2/n2469 ), .B0(\U1/aes_core/SB2/n2387 ), .Y(
        \U1/aes_core/SB2/n2202 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U790  ( .A(\U1/aes_core/SB2/n2443 ), .B(
        \U1/aes_core/SB2/n2490 ), .Y(\U1/aes_core/SB2/n2454 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U789  ( .A0(\U1/aes_core/SB2/n2308 ), 
        .A1(\U1/aes_core/SB2/n2512 ), .B0(\U1/aes_core/SB2/n2454 ), .B1(
        \U1/aes_core/SB2/n2465 ), .C0(\U1/aes_core/SB2/n2506 ), .C1(
        \U1/aes_core/SB2/n2515 ), .Y(\U1/aes_core/SB2/n2204 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U788  ( .A(\U1/aes_core/SB2/n2209 ), .B(
        \U1/aes_core/SB2/n2208 ), .C(\U1/aes_core/SB2/n2207 ), .D(
        \U1/aes_core/SB2/n2206 ), .E(\U1/aes_core/SB2/n2205 ), .F(
        \U1/aes_core/SB2/n2204 ), .Y(\U1/aes_core/SB2/n2417 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U787  ( .AN(\U1/aes_core/SB2/n2213 ), 
        .B(\U1/aes_core/SB2/n2212 ), .C(\U1/aes_core/SB2/n2211 ), .D(
        \U1/aes_core/SB2/n2210 ), .Y(\U1/aes_core/SB2/n2223 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U786  ( .A0(\U1/aes_core/SB2/n2500 ), 
        .A1(\U1/aes_core/SB2/n2410 ), .B0(\U1/aes_core/SB2/n2495 ), .B1(
        \U1/aes_core/SB2/n2409 ), .C0(\U1/aes_core/SB2/n2214 ), .C1(
        \U1/aes_core/SB2/n2510 ), .Y(\U1/aes_core/SB2/n2222 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U785  ( .A0(\U1/aes_core/SB2/n2464 ), 
        .A1(\U1/aes_core/SB2/n2370 ), .B0(\U1/aes_core/SB2/n2215 ), .B1(
        \U1/aes_core/SB2/n2308 ), .Y(\U1/aes_core/SB2/n2216 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U784  ( .A0(\U1/aes_core/SB2/n2387 ), 
        .A1(\U1/aes_core/SB2/n2404 ), .B0(\U1/aes_core/SB2/n2403 ), .B1(
        \U1/aes_core/SB2/n2467 ), .C0(\U1/aes_core/SB2/n2216 ), .Y(
        \U1/aes_core/SB2/n2221 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U783  ( .A(\U1/aes_core/SB2/n2475 ), .B(
        \U1/aes_core/SB2/n2514 ), .Y(\U1/aes_core/SB2/n2218 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U782  ( .A0(\U1/aes_core/SB2/n2300 ), 
        .A1(\U1/aes_core/SB2/n2219 ), .B0(\U1/aes_core/SB2/n2496 ), .B1(
        \U1/aes_core/SB2/n2218 ), .C0(\U1/aes_core/SB2/n2217 ), .Y(
        \U1/aes_core/SB2/n2220 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U781  ( .AN(\U1/aes_core/SB2/n2223 ), 
        .B(\U1/aes_core/SB2/n2222 ), .C(\U1/aes_core/SB2/n2221 ), .D(
        \U1/aes_core/SB2/n2220 ), .Y(\U1/aes_core/SB2/n2462 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U780  ( .A(\U1/aes_core/SB2/n2224 ), .Y(
        \U1/aes_core/SB2/n2240 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U779  ( .A0(\U1/aes_core/SB2/n2354 ), 
        .A1(\U1/aes_core/SB2/n2423 ), .B0(\U1/aes_core/SB2/n2225 ), .Y(
        \U1/aes_core/SB2/n2239 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U778  ( .A0(\U1/aes_core/SB2/n2496 ), 
        .A1(\U1/aes_core/SB2/n2495 ), .B0(\U1/aes_core/SB2/n2466 ), .B1(
        \U1/aes_core/SB2/n2226 ), .Y(\U1/aes_core/SB2/n2227 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U777  ( .A0(\U1/aes_core/SB2/n2477 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2493 ), .B1(
        \U1/aes_core/SB2/n2505 ), .C0(\U1/aes_core/SB2/n2227 ), .Y(
        \U1/aes_core/SB2/n2238 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U776  ( .A(\U1/aes_core/SB2/n2231 ), .B(
        \U1/aes_core/SB2/n2230 ), .C(\U1/aes_core/SB2/n2229 ), .D(
        \U1/aes_core/SB2/n2228 ), .Y(\U1/aes_core/SB2/n2237 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U775  ( .AN(\U1/aes_core/SB2/n2235 ), 
        .B(\U1/aes_core/SB2/n2234 ), .C(\U1/aes_core/SB2/n2233 ), .D(
        \U1/aes_core/SB2/n2232 ), .Y(\U1/aes_core/SB2/n2236 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U774  ( .A(\U1/aes_core/SB2/n2241 ), .B(
        \U1/aes_core/SB2/n2240 ), .C(\U1/aes_core/SB2/n2239 ), .D(
        \U1/aes_core/SB2/n2238 ), .E(\U1/aes_core/SB2/n2237 ), .F(
        \U1/aes_core/SB2/n2236 ), .Y(\U1/aes_core/SB2/n2366 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U773  ( .A0(\U1/aes_core/SB2/n2453 ), 
        .A1(\U1/aes_core/SB2/n2370 ), .B0(\U1/aes_core/SB2/n2242 ), .Y(
        \U1/aes_core/SB2/n2257 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U772  ( .AN(\U1/aes_core/SB2/n2246 ), 
        .B(\U1/aes_core/SB2/n2245 ), .C(\U1/aes_core/SB2/n2244 ), .D(
        \U1/aes_core/SB2/n2243 ), .Y(\U1/aes_core/SB2/n2256 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U771  ( .A(\U1/aes_core/SB2/n2487 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2501 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U770  ( .A(\U1/aes_core/SB2/n2249 ), .B(
        \U1/aes_core/SB2/n2248 ), .C(\U1/aes_core/SB2/n2247 ), .D(
        \U1/aes_core/SB2/n2501 ), .Y(\U1/aes_core/SB2/n2255 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U769  ( .A(\U1/aes_core/SB2/n2253 ), .B(
        \U1/aes_core/SB2/n2252 ), .C(\U1/aes_core/SB2/n2251 ), .D(
        \U1/aes_core/SB2/n2250 ), .Y(\U1/aes_core/SB2/n2254 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U768  ( .A(\U1/aes_core/SB2/n2259 ), .B(
        \U1/aes_core/SB2/n2258 ), .C(\U1/aes_core/SB2/n2257 ), .D(
        \U1/aes_core/SB2/n2256 ), .E(\U1/aes_core/SB2/n2255 ), .F(
        \U1/aes_core/SB2/n2254 ), .Y(\U1/aes_core/SB2/n2390 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U767  ( .AN(\U1/aes_core/SB2/n2263 ), 
        .B(\U1/aes_core/SB2/n2262 ), .C(\U1/aes_core/SB2/n2261 ), .D(
        \U1/aes_core/SB2/n2260 ), .Y(\U1/aes_core/SB2/n2272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U766  ( .A(\U1/aes_core/SB2/n2267 ), .B(
        \U1/aes_core/SB2/n2266 ), .C(\U1/aes_core/SB2/n2265 ), .D(
        \U1/aes_core/SB2/n2264 ), .Y(\U1/aes_core/SB2/n2271 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U765  ( .A(\U1/aes_core/SB2/n2452 ), .B(
        \U1/aes_core/SB2/n2488 ), .C(\U1/aes_core/SB2/n2490 ), .Y(
        \U1/aes_core/SB2/n2269 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U764  ( .A0(\U1/aes_core/SB2/n2269 ), 
        .A1(\U1/aes_core/SB2/n2478 ), .B0(\U1/aes_core/SB2/n2308 ), .B1(
        \U1/aes_core/SB2/n2514 ), .C0(\U1/aes_core/SB2/n2268 ), .Y(
        \U1/aes_core/SB2/n2270 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U763  ( .A(\U1/aes_core/SB2/n2275 ), .B(
        \U1/aes_core/SB2/n2274 ), .C(\U1/aes_core/SB2/n2273 ), .D(
        \U1/aes_core/SB2/n2272 ), .E(\U1/aes_core/SB2/n2271 ), .F(
        \U1/aes_core/SB2/n2270 ), .Y(\U1/aes_core/SB2/n2438 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U762  ( .A0(\U1/aes_core/SB2/n2308 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2276 ), .Y(
        \U1/aes_core/SB2/n2290 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U761  ( .A0(\U1/aes_core/SB2/n2442 ), 
        .A1(\U1/aes_core/SB2/n2444 ), .B0(\U1/aes_core/SB2/n2499 ), .B1(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U760  ( .A0(\U1/aes_core/SB2/n2353 ), 
        .A1(\U1/aes_core/SB2/n2441 ), .B0(\U1/aes_core/SB2/n2354 ), .B1(
        \U1/aes_core/SB2/n2418 ), .C0(\U1/aes_core/SB2/n2277 ), .Y(
        \U1/aes_core/SB2/n2289 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U759  ( .A(\U1/aes_core/SB2/n2278 ), .Y(
        \U1/aes_core/SB2/n2281 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U758  ( .AN(\U1/aes_core/SB2/n2282 ), 
        .B(\U1/aes_core/SB2/n2281 ), .C(\U1/aes_core/SB2/n2280 ), .D(
        \U1/aes_core/SB2/n2279 ), .Y(\U1/aes_core/SB2/n2288 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U757  ( .A(\U1/aes_core/SB2/n2286 ), .B(
        \U1/aes_core/SB2/n2285 ), .C(\U1/aes_core/SB2/n2284 ), .D(
        \U1/aes_core/SB2/n2283 ), .Y(\U1/aes_core/SB2/n2287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U756  ( .A(\U1/aes_core/SB2/n2292 ), .B(
        \U1/aes_core/SB2/n2291 ), .C(\U1/aes_core/SB2/n2290 ), .D(
        \U1/aes_core/SB2/n2289 ), .E(\U1/aes_core/SB2/n2288 ), .F(
        \U1/aes_core/SB2/n2287 ), .Y(\U1/aes_core/SB2/n2397 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U755  ( .A0(\U1/aes_core/SB2/n2488 ), 
        .A1(\U1/aes_core/SB2/n2293 ), .B0(\U1/aes_core/SB2/n2498 ), .B1(
        \U1/aes_core/SB2/n2444 ), .Y(\U1/aes_core/SB2/n2294 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U754  ( .A0(\U1/aes_core/SB2/n2370 ), 
        .A1(\U1/aes_core/SB2/n2515 ), .B0(\U1/aes_core/SB2/n2295 ), .B1(
        \U1/aes_core/SB2/n2505 ), .C0(\U1/aes_core/SB2/n2294 ), .Y(
        \U1/aes_core/SB2/n2307 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U753  ( .AN(\U1/aes_core/SB2/n2299 ), 
        .B(\U1/aes_core/SB2/n2298 ), .C(\U1/aes_core/SB2/n2297 ), .D(
        \U1/aes_core/SB2/n2296 ), .Y(\U1/aes_core/SB2/n2306 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U752  ( .A0(\U1/aes_core/SB2/n2508 ), 
        .A1(\U1/aes_core/SB2/n2300 ), .B0(\U1/aes_core/SB2/n2499 ), .Y(
        \U1/aes_core/SB2/n2304 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U751  ( .A(\U1/aes_core/SB2/n2475 ), .B(
        \U1/aes_core/SB2/n2480 ), .Y(\U1/aes_core/SB2/n2301 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U750  ( .A0(\U1/aes_core/SB2/n2451 ), 
        .A1(\U1/aes_core/SB2/n2301 ), .B0(\U1/aes_core/SB2/n2452 ), .B1(
        \U1/aes_core/SB2/n2398 ), .Y(\U1/aes_core/SB2/n2302 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U749  ( .A(\U1/aes_core/SB2/n2304 ), .B(
        \U1/aes_core/SB2/n2303 ), .C(\U1/aes_core/SB2/n2302 ), .Y(
        \U1/aes_core/SB2/n2305 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U748  ( .A(\U1/aes_core/SB2/n2390 ), .B(
        \U1/aes_core/SB2/n2438 ), .C(\U1/aes_core/SB2/n2397 ), .D(
        \U1/aes_core/SB2/n2307 ), .E(\U1/aes_core/SB2/n2306 ), .F(
        \U1/aes_core/SB2/n2305 ), .Y(\U1/aes_core/SB2/n2484 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U747  ( .A(\U1/aes_core/SB2/n2417 ), .B(
        \U1/aes_core/SB2/n2462 ), .C(\U1/aes_core/SB2/n2366 ), .D(
        \U1/aes_core/SB2/n2484 ), .Y(\U1/aes_core/SB2/n2321 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U746  ( .A0(\U1/aes_core/SB2/n2464 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2308 ), .B1(
        \U1/aes_core/SB2/n2480 ), .Y(\U1/aes_core/SB2/n2309 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U745  ( .A0(\U1/aes_core/SB2/n2469 ), 
        .A1(\U1/aes_core/SB2/n2487 ), .B0(\U1/aes_core/SB2/n2500 ), .B1(
        \U1/aes_core/SB2/n2508 ), .C0(\U1/aes_core/SB2/n2309 ), .Y(
        \U1/aes_core/SB2/n2320 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U744  ( .A(\U1/aes_core/SB2/n2310 ), .Y(
        \U1/aes_core/SB2/n2313 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U743  ( .A0(\U1/aes_core/SB2/n2311 ), 
        .A1(\U1/aes_core/SB2/n2441 ), .B0(\U1/aes_core/SB2/n2369 ), .B1(
        \U1/aes_core/SB2/n2421 ), .Y(\U1/aes_core/SB2/n2312 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U742  ( .A0(\U1/aes_core/SB2/n2488 ), 
        .A1(\U1/aes_core/SB2/n2313 ), .B0(\U1/aes_core/SB2/n2470 ), .B1(
        \U1/aes_core/SB2/n2419 ), .C0(\U1/aes_core/SB2/n2312 ), .Y(
        \U1/aes_core/SB2/n2319 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U741  ( .A0(\U1/aes_core/SB2/n2510 ), 
        .A1(\U1/aes_core/SB2/n2387 ), .B0(\U1/aes_core/SB2/n2490 ), .Y(
        \U1/aes_core/SB2/n2317 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB2/U740  ( .A(\U1/aes_core/SB2/n2317 ), .B(
        \U1/aes_core/SB2/n2316 ), .C(\U1/aes_core/SB2/n2315 ), .D(
        \U1/aes_core/SB2/n2314 ), .Y(\U1/aes_core/SB2/n2318 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U739  ( .AN(\U1/aes_core/SB2/n2321 ), 
        .B(\U1/aes_core/SB2/n2320 ), .C(\U1/aes_core/SB2/n2319 ), .D(
        \U1/aes_core/SB2/n2318 ), .Y(\U1/aes_core/sb2 [19]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U738  ( .A(\U1/aes_core/SB2/n3166 ), .B(
        \U1/aes_core/SB2/n2983 ), .Y(\U1/aes_core/SB2/n3043 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U737  ( .A(\U1/aes_core/SB2/n3113 ), .B(
        \U1/aes_core/SB2/n3163 ), .Y(\U1/aes_core/SB2/n3003 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U736  ( .A(\U1/aes_core/SB2/n3130 ), .B(
        \U1/aes_core/SB2/n3241 ), .Y(\U1/aes_core/SB2/n3112 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U735  ( .A0(\U1/aes_core/SB2/n3112 ), 
        .A1(\U1/aes_core/SB2/n3166 ), .B0(\U1/aes_core/SB2/n3255 ), .Y(
        \U1/aes_core/SB2/n2326 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U734  ( .A(\U1/aes_core/SB2/n3194 ), .B(
        \U1/aes_core/SB2/n3242 ), .Y(\U1/aes_core/SB2/n3019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U733  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3194 ), .Y(\U1/aes_core/SB2/n3118 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U732  ( .A(\U1/aes_core/SB2/n3239 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3051 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U731  ( .A(\U1/aes_core/SB2/n3019 ), .B(
        \U1/aes_core/SB2/n3118 ), .C(\U1/aes_core/SB2/n3051 ), .Y(
        \U1/aes_core/SB2/n2325 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U730  ( .A(\U1/aes_core/SB2/n3194 ), .B(
        \U1/aes_core/SB2/n3253 ), .Y(\U1/aes_core/SB2/n3078 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U729  ( .A(\U1/aes_core/SB2/n3239 ), .B(
        \U1/aes_core/SB2/n3230 ), .C(\U1/aes_core/SB2/n3251 ), .Y(
        \U1/aes_core/SB2/n2322 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U728  ( .A0(\U1/aes_core/SB2/n3078 ), 
        .A1(\U1/aes_core/SB2/n3219 ), .B0(\U1/aes_core/SB2/n2322 ), .B1(
        \U1/aes_core/SB2/n3249 ), .C0(\U1/aes_core/SB2/n3113 ), .C1(
        \U1/aes_core/SB2/n3145 ), .Y(\U1/aes_core/SB2/n2324 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U727  ( .A0(\U1/aes_core/SB2/n3220 ), 
        .A1(\U1/aes_core/SB2/n3248 ), .B0(\U1/aes_core/SB2/n3221 ), .B1(
        \U1/aes_core/SB2/n3218 ), .Y(\U1/aes_core/SB2/n2323 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U726  ( .A(\U1/aes_core/SB2/n3043 ), .B(
        \U1/aes_core/SB2/n3003 ), .C(\U1/aes_core/SB2/n2326 ), .D(
        \U1/aes_core/SB2/n2325 ), .E(\U1/aes_core/SB2/n2324 ), .F(
        \U1/aes_core/SB2/n2323 ), .Y(\U1/aes_core/SB2/n3263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U725  ( .A(\U1/aes_core/SB2/n3094 ), .B(
        \U1/aes_core/SB2/n3079 ), .Y(\U1/aes_core/SB2/n2969 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U724  ( .A0(\U1/aes_core/SB2/n3094 ), 
        .A1(\U1/aes_core/SB2/n3184 ), .B0(\U1/aes_core/SB2/n2983 ), .Y(
        \U1/aes_core/SB2/n2333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U723  ( .A(\U1/aes_core/SB2/n3188 ), .B(
        \U1/aes_core/SB2/n3194 ), .Y(\U1/aes_core/SB2/n2971 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U722  ( .A0(\U1/aes_core/SB2/n3076 ), 
        .A1(\U1/aes_core/SB2/n3223 ), .B0(\U1/aes_core/SB2/n2971 ), .B1(
        \U1/aes_core/SB2/n3237 ), .Y(\U1/aes_core/SB2/n2332 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U721  ( .A0(\U1/aes_core/SB2/n3063 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3207 ), .B1(
        \U1/aes_core/SB2/n3113 ), .C0(\U1/aes_core/SB2/n3221 ), .C1(
        \U1/aes_core/SB2/n3164 ), .Y(\U1/aes_core/SB2/n2331 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U720  ( .A(\U1/aes_core/SB2/n3256 ), .B(
        \U1/aes_core/SB2/n2327 ), .Y(\U1/aes_core/SB2/n3027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U719  ( .A(\U1/aes_core/SB2/n3243 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U718  ( .A(\U1/aes_core/SB2/n3185 ), .B(
        \U1/aes_core/SB2/n3238 ), .Y(\U1/aes_core/SB2/n3044 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U717  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3253 ), .Y(\U1/aes_core/SB2/n3148 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U716  ( .AN(\U1/aes_core/SB2/n3027 ), 
        .B(\U1/aes_core/SB2/n3034 ), .C(\U1/aes_core/SB2/n3044 ), .D(
        \U1/aes_core/SB2/n3148 ), .Y(\U1/aes_core/SB2/n2330 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U715  ( .A(\U1/aes_core/SB2/n3145 ), .B(
        \U1/aes_core/SB2/n2328 ), .Y(\U1/aes_core/SB2/n3127 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U714  ( .A(\U1/aes_core/SB2/n3223 ), .B(
        \U1/aes_core/SB2/n3207 ), .Y(\U1/aes_core/SB2/n3180 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U712  ( .A(\U1/aes_core/SB2/n2968 ), .B(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n2993 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U710  ( .A(\U1/aes_core/SB2/n2969 ), .B(
        \U1/aes_core/SB2/n2333 ), .C(\U1/aes_core/SB2/n2332 ), .D(
        \U1/aes_core/SB2/n2331 ), .E(\U1/aes_core/SB2/n2330 ), .F(
        \U1/aes_core/SB2/n2329 ), .Y(\U1/aes_core/SB2/n2904 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U709  ( .A(\U1/aes_core/SB2/n3161 ), .B(
        \U1/aes_core/SB2/n2983 ), .Y(\U1/aes_core/SB2/n2981 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U708  ( .A(\U1/aes_core/SB2/n3113 ), .B(
        \U1/aes_core/SB2/n3063 ), .Y(\U1/aes_core/SB2/n3193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U707  ( .A(\U1/aes_core/SB2/n3094 ), .B(
        \U1/aes_core/SB2/n3164 ), .Y(\U1/aes_core/SB2/n3031 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U706  ( .A(\U1/aes_core/SB2/n3258 ), .B(
        \U1/aes_core/SB2/n3164 ), .Y(\U1/aes_core/SB2/n3046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U705  ( .A(\U1/aes_core/SB2/n3189 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n3106 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U704  ( .A(\U1/aes_core/SB2/n3239 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n2998 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U703  ( .A(\U1/aes_core/SB2/n3243 ), .B(
        \U1/aes_core/SB2/n3239 ), .Y(\U1/aes_core/SB2/n3092 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U702  ( .A(\U1/aes_core/SB2/n3153 ), .B(
        \U1/aes_core/SB2/n3210 ), .Y(\U1/aes_core/SB2/n3017 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U701  ( .A(\U1/aes_core/SB2/n3106 ), .B(
        \U1/aes_core/SB2/n2998 ), .C(\U1/aes_core/SB2/n3092 ), .D(
        \U1/aes_core/SB2/n3017 ), .Y(\U1/aes_core/SB2/n2337 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U700  ( .A(\U1/aes_core/SB2/n3258 ), .B(
        \U1/aes_core/SB2/n3079 ), .Y(\U1/aes_core/SB2/n3067 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U699  ( .A(\U1/aes_core/SB2/n3257 ), .B(
        \U1/aes_core/SB2/n3063 ), .Y(\U1/aes_core/SB2/n3167 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U698  ( .A(\U1/aes_core/SB2/n3184 ), .B(
        \U1/aes_core/SB2/n3223 ), .Y(\U1/aes_core/SB2/n3117 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U697  ( .A(\U1/aes_core/SB2/n3145 ), .B(
        \U1/aes_core/SB2/n3223 ), .Y(\U1/aes_core/SB2/n2967 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U696  ( .A0(\U1/aes_core/SB2/n3223 ), 
        .A1(\U1/aes_core/SB2/n3258 ), .B0(\U1/aes_core/SB2/n3079 ), .B1(
        \U1/aes_core/SB2/n3184 ), .Y(\U1/aes_core/SB2/n2335 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U695  ( .A0(\U1/aes_core/SB2/n3063 ), 
        .A1(\U1/aes_core/SB2/n3255 ), .B0(\U1/aes_core/SB2/n3076 ), .B1(
        \U1/aes_core/SB2/n3113 ), .Y(\U1/aes_core/SB2/n2334 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U694  ( .A(\U1/aes_core/SB2/n3067 ), .B(
        \U1/aes_core/SB2/n3167 ), .C(\U1/aes_core/SB2/n3117 ), .D(
        \U1/aes_core/SB2/n2967 ), .E(\U1/aes_core/SB2/n2335 ), .F(
        \U1/aes_core/SB2/n2334 ), .Y(\U1/aes_core/SB2/n2336 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U693  ( .A(\U1/aes_core/SB2/n2981 ), .B(
        \U1/aes_core/SB2/n3193 ), .C(\U1/aes_core/SB2/n3031 ), .D(
        \U1/aes_core/SB2/n3046 ), .E(\U1/aes_core/SB2/n2337 ), .F(
        \U1/aes_core/SB2/n2336 ), .Y(\U1/aes_core/SB2/n2893 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U692  ( .A0(\U1/aes_core/SB2/n3189 ), 
        .A1(\U1/aes_core/SB2/n3186 ), .B0(\U1/aes_core/SB2/n3242 ), .B1(
        \U1/aes_core/SB2/n3130 ), .C0(\U1/aes_core/SB2/n2893 ), .Y(
        \U1/aes_core/SB2/n2338 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U691  ( .A(\U1/aes_core/SB2/n2338 ), .Y(
        \U1/aes_core/SB2/n2345 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U690  ( .A(\U1/aes_core/SB2/n3221 ), .B(
        \U1/aes_core/SB2/n3184 ), .Y(\U1/aes_core/SB2/n3211 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U689  ( .A0(\U1/aes_core/SB2/n3188 ), 
        .A1(\U1/aes_core/SB2/n3211 ), .B0(\U1/aes_core/SB2/n3243 ), .Y(
        \U1/aes_core/SB2/n2341 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U688  ( .A0(\U1/aes_core/SB2/n3153 ), 
        .A1(\U1/aes_core/SB2/n3232 ), .B0(\U1/aes_core/SB2/n3195 ), .Y(
        \U1/aes_core/SB2/n2340 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U687  ( .A0(\U1/aes_core/SB2/n3152 ), 
        .A1(\U1/aes_core/SB2/n3194 ), .B0(\U1/aes_core/SB2/n3238 ), .Y(
        \U1/aes_core/SB2/n2339 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U686  ( .A(\U1/aes_core/SB2/n3185 ), .B(
        \U1/aes_core/SB2/n3231 ), .Y(\U1/aes_core/SB2/n3010 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U685  ( .A(\U1/aes_core/SB2/n2341 ), .B(
        \U1/aes_core/SB2/n2340 ), .C(\U1/aes_core/SB2/n2339 ), .D(
        \U1/aes_core/SB2/n3010 ), .Y(\U1/aes_core/SB2/n2344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U684  ( .A(\U1/aes_core/SB2/n3230 ), .B(
        \U1/aes_core/SB2/n3146 ), .Y(\U1/aes_core/SB2/n3200 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB2/U683  ( .A(\U1/aes_core/SB2/n3200 ), .B(
        \U1/aes_core/SB2/n3220 ), .C(\U1/aes_core/SB2/n3207 ), .Y(
        \U1/aes_core/SB2/n2342 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U682  ( .A0(\U1/aes_core/SB2/n3184 ), 
        .A1(\U1/aes_core/SB2/n3257 ), .B0(\U1/aes_core/SB2/n2342 ), .B1(
        \U1/aes_core/SB2/n3218 ), .C0(\U1/aes_core/SB2/n3256 ), .C1(
        \U1/aes_core/SB2/n3248 ), .Y(\U1/aes_core/SB2/n2343 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U681  ( .A(\U1/aes_core/SB2/n3263 ), .B(
        \U1/aes_core/SB2/n2904 ), .C(\U1/aes_core/SB2/n2346 ), .D(
        \U1/aes_core/SB2/n2345 ), .E(\U1/aes_core/SB2/n2344 ), .F(
        \U1/aes_core/SB2/n2343 ), .Y(\U1/aes_core/sb2 [1]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U680  ( .A0(\U1/aes_core/SB2/n2361 ), 
        .A1(\U1/aes_core/SB2/n2476 ), .B0(\U1/aes_core/SB2/n2420 ), .Y(
        \U1/aes_core/SB2/n2358 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U679  ( .A(\U1/aes_core/SB2/n2349 ), .B(
        \U1/aes_core/SB2/n2348 ), .C(\U1/aes_core/SB2/n2347 ), .Y(
        \U1/aes_core/SB2/n2357 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U678  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2499 ), .Y(\U1/aes_core/SB2/n2352 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U677  ( .A(\U1/aes_core/SB2/n2470 ), .B(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2350 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U676  ( .A0(\U1/aes_core/SB2/n2352 ), 
        .A1(\U1/aes_core/SB2/n2351 ), .B0(\U1/aes_core/SB2/n2350 ), .B1(
        \U1/aes_core/SB2/n2493 ), .C0(\U1/aes_core/SB2/n2476 ), .C1(
        \U1/aes_core/SB2/n2402 ), .Y(\U1/aes_core/SB2/n2356 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U675  ( .A0(\U1/aes_core/SB2/n2453 ), 
        .A1(\U1/aes_core/SB2/n2354 ), .B0(\U1/aes_core/SB2/n2515 ), .B1(
        \U1/aes_core/SB2/n2505 ), .C0(\U1/aes_core/SB2/n2478 ), .C1(
        \U1/aes_core/SB2/n2353 ), .Y(\U1/aes_core/SB2/n2355 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U674  ( .A(\U1/aes_core/SB2/n2360 ), .B(
        \U1/aes_core/SB2/n2359 ), .C(\U1/aes_core/SB2/n2358 ), .D(
        \U1/aes_core/SB2/n2357 ), .E(\U1/aes_core/SB2/n2356 ), .F(
        \U1/aes_core/SB2/n2355 ), .Y(\U1/aes_core/SB2/n2485 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U673  ( .A0(\U1/aes_core/SB2/n2361 ), 
        .A1(\U1/aes_core/SB2/n2370 ), .B0(\U1/aes_core/SB2/n2441 ), .Y(
        \U1/aes_core/SB2/n2396 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB2/U672  ( .A0(\U1/aes_core/SB2/n2465 ), 
        .A1(\U1/aes_core/SB2/n2478 ), .A2(\U1/aes_core/SB2/n2418 ), .B0(
        \U1/aes_core/SB2/n2494 ), .Y(\U1/aes_core/SB2/n2395 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U671  ( .A(\U1/aes_core/SB2/n2365 ), .B(
        \U1/aes_core/SB2/n2364 ), .C(\U1/aes_core/SB2/n2363 ), .D(
        \U1/aes_core/SB2/n2362 ), .Y(\U1/aes_core/SB2/n2392 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U670  ( .A(\U1/aes_core/SB2/n2366 ), .Y(
        \U1/aes_core/SB2/n2389 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U669  ( .A(\U1/aes_core/SB2/n2367 ), .Y(
        \U1/aes_core/SB2/n2383 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB2/U668  ( .A0(\U1/aes_core/SB2/n2369 ), 
        .A1(\U1/aes_core/SB2/n2506 ), .B0N(\U1/aes_core/SB2/n2368 ), .Y(
        \U1/aes_core/SB2/n2382 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U667  ( .A0(\U1/aes_core/SB2/n2513 ), 
        .A1(\U1/aes_core/SB2/n2370 ), .B0(\U1/aes_core/SB2/n2420 ), .B1(
        \U1/aes_core/SB2/n2480 ), .C0(\U1/aes_core/SB2/n2494 ), .C1(
        \U1/aes_core/SB2/n2515 ), .Y(\U1/aes_core/SB2/n2381 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U666  ( .AN(\U1/aes_core/SB2/n2374 ), 
        .B(\U1/aes_core/SB2/n2373 ), .C(\U1/aes_core/SB2/n2372 ), .D(
        \U1/aes_core/SB2/n2371 ), .Y(\U1/aes_core/SB2/n2380 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U665  ( .A(\U1/aes_core/SB2/n2378 ), .B(
        \U1/aes_core/SB2/n2377 ), .C(\U1/aes_core/SB2/n2376 ), .D(
        \U1/aes_core/SB2/n2375 ), .Y(\U1/aes_core/SB2/n2379 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U664  ( .A(\U1/aes_core/SB2/n2384 ), .B(
        \U1/aes_core/SB2/n2383 ), .C(\U1/aes_core/SB2/n2382 ), .D(
        \U1/aes_core/SB2/n2381 ), .E(\U1/aes_core/SB2/n2380 ), .F(
        \U1/aes_core/SB2/n2379 ), .Y(\U1/aes_core/SB2/n2385 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U663  ( .A(\U1/aes_core/SB2/n2385 ), .Y(
        \U1/aes_core/SB2/n2463 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U662  ( .A0(\U1/aes_core/SB2/n2453 ), 
        .A1(\U1/aes_core/SB2/n2475 ), .B0(\U1/aes_core/SB2/n2515 ), .B1(
        \U1/aes_core/SB2/n2514 ), .Y(\U1/aes_core/SB2/n2386 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U661  ( .A0(\U1/aes_core/SB2/n2443 ), 
        .A1(\U1/aes_core/SB2/n2387 ), .B0(\U1/aes_core/SB2/n2467 ), .B1(
        \U1/aes_core/SB2/n2489 ), .C0(\U1/aes_core/SB2/n2386 ), .Y(
        \U1/aes_core/SB2/n2388 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U660  ( .AN(\U1/aes_core/SB2/n2390 ), 
        .B(\U1/aes_core/SB2/n2389 ), .C(\U1/aes_core/SB2/n2463 ), .D(
        \U1/aes_core/SB2/n2388 ), .Y(\U1/aes_core/SB2/n2391 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U659  ( .A(\U1/aes_core/SB2/n2396 ), .B(
        \U1/aes_core/SB2/n2395 ), .C(\U1/aes_core/SB2/n2394 ), .D(
        \U1/aes_core/SB2/n2393 ), .E(\U1/aes_core/SB2/n2392 ), .F(
        \U1/aes_core/SB2/n2391 ), .Y(\U1/aes_core/SB2/n2461 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U658  ( .A(\U1/aes_core/SB2/n2397 ), .Y(
        \U1/aes_core/SB2/n2401 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U657  ( .A0(\U1/aes_core/SB2/n2399 ), 
        .A1(\U1/aes_core/SB2/n2398 ), .B0(\U1/aes_core/SB2/n2445 ), .B1(
        \U1/aes_core/SB2/n2404 ), .Y(\U1/aes_core/SB2/n2400 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U656  ( .A0(\U1/aes_core/SB2/n2494 ), 
        .A1(\U1/aes_core/SB2/n2402 ), .B0(\U1/aes_core/SB2/n2401 ), .C0(
        \U1/aes_core/SB2/n2400 ), .Y(\U1/aes_core/SB2/n2416 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U655  ( .A0(\U1/aes_core/SB2/n2403 ), 
        .A1(\U1/aes_core/SB2/n2466 ), .B0(\U1/aes_core/SB2/n2495 ), .Y(
        \U1/aes_core/SB2/n2408 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U654  ( .A0(\U1/aes_core/SB2/n2404 ), 
        .A1(\U1/aes_core/SB2/n2469 ), .B0(\U1/aes_core/SB2/n2498 ), .Y(
        \U1/aes_core/SB2/n2407 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U653  ( .A(\U1/aes_core/SB2/n2408 ), .B(
        \U1/aes_core/SB2/n2407 ), .C(\U1/aes_core/SB2/n2406 ), .D(
        \U1/aes_core/SB2/n2405 ), .Y(\U1/aes_core/SB2/n2415 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U652  ( .A(\U1/aes_core/SB2/n2446 ), .B(
        \U1/aes_core/SB2/n2409 ), .Y(\U1/aes_core/SB2/n2413 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U651  ( .A(\U1/aes_core/SB2/n2410 ), .B(
        \U1/aes_core/SB2/n2451 ), .Y(\U1/aes_core/SB2/n2412 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U650  ( .A0(\U1/aes_core/SB2/n2413 ), 
        .A1(\U1/aes_core/SB2/n2512 ), .B0(\U1/aes_core/SB2/n2412 ), .B1(
        \U1/aes_core/SB2/n2476 ), .C0(\U1/aes_core/SB2/n2411 ), .C1(
        \U1/aes_core/SB2/n2477 ), .Y(\U1/aes_core/SB2/n2414 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U649  ( .A(\U1/aes_core/SB2/n2485 ), .B(
        \U1/aes_core/SB2/n2461 ), .C(\U1/aes_core/SB2/n2417 ), .D(
        \U1/aes_core/SB2/n2416 ), .E(\U1/aes_core/SB2/n2415 ), .F(
        \U1/aes_core/SB2/n2414 ), .Y(\U1/aes_core/sb2 [20]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U648  ( .A1N(\U1/aes_core/SB2/n2419 ), 
        .A0(\U1/aes_core/SB2/n2418 ), .B0(\U1/aes_core/SB2/n2475 ), .Y(
        \U1/aes_core/SB2/n2435 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U647  ( .A(\U1/aes_core/SB2/n2488 ), .B(
        \U1/aes_core/SB2/n2469 ), .Y(\U1/aes_core/SB2/n2422 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U646  ( .A0(\U1/aes_core/SB2/n2512 ), 
        .A1(\U1/aes_core/SB2/n2423 ), .B0(\U1/aes_core/SB2/n2422 ), .B1(
        \U1/aes_core/SB2/n2515 ), .C0(\U1/aes_core/SB2/n2421 ), .C1(
        \U1/aes_core/SB2/n2420 ), .Y(\U1/aes_core/SB2/n2434 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U645  ( .A(\U1/aes_core/SB2/n2424 ), .Y(
        \U1/aes_core/SB2/n2427 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U644  ( .AN(\U1/aes_core/SB2/n2428 ), 
        .B(\U1/aes_core/SB2/n2427 ), .C(\U1/aes_core/SB2/n2426 ), .D(
        \U1/aes_core/SB2/n2425 ), .Y(\U1/aes_core/SB2/n2433 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U643  ( .A(\U1/aes_core/SB2/n2431 ), .B(
        \U1/aes_core/SB2/n2430 ), .C(\U1/aes_core/SB2/n2429 ), .Y(
        \U1/aes_core/SB2/n2432 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U642  ( .A(\U1/aes_core/SB2/n2437 ), .B(
        \U1/aes_core/SB2/n2436 ), .C(\U1/aes_core/SB2/n2435 ), .D(
        \U1/aes_core/SB2/n2434 ), .E(\U1/aes_core/SB2/n2433 ), .F(
        \U1/aes_core/SB2/n2432 ), .Y(\U1/aes_core/SB2/n2486 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U641  ( .A(\U1/aes_core/SB2/n2438 ), .Y(
        \U1/aes_core/SB2/n2440 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U640  ( .A0(\U1/aes_core/SB2/n2499 ), 
        .A1(\U1/aes_core/SB2/n2496 ), .B0(\U1/aes_core/SB2/n2500 ), .B1(
        \U1/aes_core/SB2/n2498 ), .Y(\U1/aes_core/SB2/n2439 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U639  ( .A0(\U1/aes_core/SB2/n2475 ), 
        .A1(\U1/aes_core/SB2/n2441 ), .B0(\U1/aes_core/SB2/n2440 ), .C0(
        \U1/aes_core/SB2/n2439 ), .Y(\U1/aes_core/SB2/n2460 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U638  ( .A0(\U1/aes_core/SB2/n2443 ), 
        .A1(\U1/aes_core/SB2/n2499 ), .B0(\U1/aes_core/SB2/n2442 ), .Y(
        \U1/aes_core/SB2/n2449 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U637  ( .A0(\U1/aes_core/SB2/n2446 ), 
        .A1(\U1/aes_core/SB2/n2445 ), .B0(\U1/aes_core/SB2/n2444 ), .Y(
        \U1/aes_core/SB2/n2448 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U636  ( .AN(\U1/aes_core/SB2/n2450 ), 
        .B(\U1/aes_core/SB2/n2449 ), .C(\U1/aes_core/SB2/n2448 ), .D(
        \U1/aes_core/SB2/n2447 ), .Y(\U1/aes_core/SB2/n2459 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U635  ( .A0(\U1/aes_core/SB2/n2495 ), 
        .A1(\U1/aes_core/SB2/n2452 ), .B0(\U1/aes_core/SB2/n2451 ), .Y(
        \U1/aes_core/SB2/n2456 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB2/U634  ( .A0(\U1/aes_core/SB2/n2477 ), .A1(
        \U1/aes_core/SB2/n2454 ), .B0(\U1/aes_core/SB2/n2514 ), .B1(
        \U1/aes_core/SB2/n2453 ), .Y(\U1/aes_core/SB2/n2455 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U633  ( .A0(\U1/aes_core/SB2/n2457 ), 
        .A1(\U1/aes_core/SB2/n2476 ), .B0(\U1/aes_core/SB2/n2456 ), .C0(
        \U1/aes_core/SB2/n2455 ), .Y(\U1/aes_core/SB2/n2458 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U632  ( .A(\U1/aes_core/SB2/n2486 ), .B(
        \U1/aes_core/SB2/n2462 ), .C(\U1/aes_core/SB2/n2461 ), .D(
        \U1/aes_core/SB2/n2460 ), .E(\U1/aes_core/SB2/n2459 ), .F(
        \U1/aes_core/SB2/n2458 ), .Y(\U1/aes_core/sb2 [21]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U631  ( .A0(\U1/aes_core/SB2/n2465 ), 
        .A1(\U1/aes_core/SB2/n2505 ), .B0(\U1/aes_core/SB2/n2464 ), .B1(
        \U1/aes_core/SB2/n2512 ), .C0(\U1/aes_core/SB2/n2463 ), .Y(
        \U1/aes_core/SB2/n2483 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U630  ( .A0(\U1/aes_core/SB2/n2466 ), 
        .A1(\U1/aes_core/SB2/n2510 ), .B0(\U1/aes_core/SB2/n2499 ), .Y(
        \U1/aes_core/SB2/n2474 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U629  ( .A0(\U1/aes_core/SB2/n2490 ), 
        .A1(\U1/aes_core/SB2/n2467 ), .B0(\U1/aes_core/SB2/n2498 ), .Y(
        \U1/aes_core/SB2/n2473 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U628  ( .A0(\U1/aes_core/SB2/n2470 ), 
        .A1(\U1/aes_core/SB2/n2469 ), .B0(\U1/aes_core/SB2/n2468 ), .Y(
        \U1/aes_core/SB2/n2472 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U627  ( .A(\U1/aes_core/SB2/n2474 ), .B(
        \U1/aes_core/SB2/n2473 ), .C(\U1/aes_core/SB2/n2472 ), .D(
        \U1/aes_core/SB2/n2471 ), .Y(\U1/aes_core/SB2/n2482 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U626  ( .A(\U1/aes_core/SB2/n2505 ), .B(
        \U1/aes_core/SB2/n2475 ), .Y(\U1/aes_core/SB2/n2507 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U625  ( .A(\U1/aes_core/SB2/n2495 ), .B(
        \U1/aes_core/SB2/n2507 ), .Y(\U1/aes_core/SB2/n2479 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U624  ( .A0(\U1/aes_core/SB2/n2493 ), 
        .A1(\U1/aes_core/SB2/n2480 ), .B0(\U1/aes_core/SB2/n2479 ), .B1(
        \U1/aes_core/SB2/n2478 ), .C0(\U1/aes_core/SB2/n2477 ), .C1(
        \U1/aes_core/SB2/n2476 ), .Y(\U1/aes_core/SB2/n2481 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U623  ( .A(\U1/aes_core/SB2/n2486 ), .B(
        \U1/aes_core/SB2/n2485 ), .C(\U1/aes_core/SB2/n2484 ), .D(
        \U1/aes_core/SB2/n2483 ), .E(\U1/aes_core/SB2/n2482 ), .F(
        \U1/aes_core/SB2/n2481 ), .Y(\U1/aes_core/sb2 [22]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U622  ( .A0(\U1/aes_core/SB2/n2490 ), 
        .A1(\U1/aes_core/SB2/n2489 ), .B0(\U1/aes_core/SB2/n2488 ), .B1(
        \U1/aes_core/SB2/n2487 ), .Y(\U1/aes_core/SB2/n2491 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U621  ( .A0(\U1/aes_core/SB2/n2494 ), 
        .A1(\U1/aes_core/SB2/n2493 ), .B0(\U1/aes_core/SB2/n2492 ), .C0(
        \U1/aes_core/SB2/n2491 ), .Y(\U1/aes_core/SB2/n2518 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U620  ( .A1N(\U1/aes_core/SB2/n2497 ), 
        .A0(\U1/aes_core/SB2/n2496 ), .B0(\U1/aes_core/SB2/n2495 ), .Y(
        \U1/aes_core/SB2/n2504 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U619  ( .A0(\U1/aes_core/SB2/n2500 ), 
        .A1(\U1/aes_core/SB2/n2499 ), .B0(\U1/aes_core/SB2/n2498 ), .Y(
        \U1/aes_core/SB2/n2503 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U618  ( .A(\U1/aes_core/SB2/n2504 ), .B(
        \U1/aes_core/SB2/n2503 ), .C(\U1/aes_core/SB2/n2502 ), .D(
        \U1/aes_core/SB2/n2501 ), .Y(\U1/aes_core/SB2/n2517 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U617  ( .A(\U1/aes_core/SB2/n2506 ), .B(
        \U1/aes_core/SB2/n2505 ), .Y(\U1/aes_core/SB2/n2509 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U616  ( .A0(\U1/aes_core/SB2/n2510 ), 
        .A1(\U1/aes_core/SB2/n2509 ), .B0(\U1/aes_core/SB2/n2508 ), .B1(
        \U1/aes_core/SB2/n2507 ), .Y(\U1/aes_core/SB2/n2511 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U615  ( .A0(\U1/aes_core/SB2/n2515 ), 
        .A1(\U1/aes_core/SB2/n2514 ), .B0(\U1/aes_core/SB2/n2513 ), .B1(
        \U1/aes_core/SB2/n2512 ), .C0(\U1/aes_core/SB2/n2511 ), .Y(
        \U1/aes_core/SB2/n2516 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U614  ( .A(\U1/aes_core/SB2/n2521 ), .B(
        \U1/aes_core/SB2/n2520 ), .C(\U1/aes_core/SB2/n2519 ), .D(
        \U1/aes_core/SB2/n2518 ), .E(\U1/aes_core/SB2/n2517 ), .F(
        \U1/aes_core/SB2/n2516 ), .Y(\U1/aes_core/sb2 [23]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U613  ( .A(Dout[63]), .B(Dout[62]), .Y(
        \U1/aes_core/SB2/n2540 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U612  ( .A(Dout[61]), .B(Dout[60]), .Y(
        \U1/aes_core/SB2/n2531 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U611  ( .A(\U1/aes_core/SB2/n2540 ), .B(
        \U1/aes_core/SB2/n2531 ), .Y(\U1/aes_core/SB2/n2604 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U610  ( .A(Dout[57]), .Y(
        \U1/aes_core/SB2/n2525 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U609  ( .A(Dout[56]), .Y(
        \U1/aes_core/SB2/n2522 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U608  ( .A(\U1/aes_core/SB2/n2525 ), .B(
        \U1/aes_core/SB2/n2522 ), .Y(\U1/aes_core/SB2/n2532 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U607  ( .A(Dout[59]), .B(Dout[58]), .Y(
        \U1/aes_core/SB2/n2552 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U606  ( .A(\U1/aes_core/SB2/n2532 ), .B(
        \U1/aes_core/SB2/n2552 ), .Y(\U1/aes_core/SB2/n2907 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U605  ( .A(\U1/aes_core/SB2/n2604 ), .B(
        \U1/aes_core/SB2/n2907 ), .Y(\U1/aes_core/SB2/n2693 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U604  ( .A(Dout[58]), .B(Dout[59]), .Y(
        \U1/aes_core/SB2/n2535 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U603  ( .A(\U1/aes_core/SB2/n2535 ), .B(
        \U1/aes_core/SB2/n2532 ), .Y(\U1/aes_core/SB2/n2824 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U602  ( .A(Dout[63]), .Y(
        \U1/aes_core/SB2/n2528 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U601  ( .A(\U1/aes_core/SB2/n2528 ), .B(
        Dout[62]), .Y(\U1/aes_core/SB2/n2558 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U600  ( .A(\U1/aes_core/SB2/n2558 ), .B(
        \U1/aes_core/SB2/n2531 ), .Y(\U1/aes_core/SB2/n2603 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U599  ( .A(\U1/aes_core/SB2/n2824 ), .B(
        \U1/aes_core/SB2/n2603 ), .Y(\U1/aes_core/SB2/n2790 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U598  ( .A(Dout[59]), .Y(
        \U1/aes_core/SB2/n2523 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB2/U597  ( .A(Dout[58]), .B(
        \U1/aes_core/SB2/n2523 ), .Y(\U1/aes_core/SB2/n2533 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U596  ( .A(\U1/aes_core/SB2/n2532 ), .B(
        \U1/aes_core/SB2/n2533 ), .Y(\U1/aes_core/SB2/n2755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U595  ( .A(\U1/aes_core/SB2/n2755 ), .Y(
        \U1/aes_core/SB2/n2941 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U594  ( .A(Dout[60]), .Y(
        \U1/aes_core/SB2/n2524 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U593  ( .A(\U1/aes_core/SB2/n2524 ), .B(
        Dout[61]), .Y(\U1/aes_core/SB2/n2539 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U592  ( .A(Dout[62]), .Y(
        \U1/aes_core/SB2/n2527 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U591  ( .A(\U1/aes_core/SB2/n2527 ), .B(
        Dout[63]), .Y(\U1/aes_core/SB2/n2549 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U590  ( .A(\U1/aes_core/SB2/n2539 ), .B(
        \U1/aes_core/SB2/n2549 ), .Y(\U1/aes_core/SB2/n2776 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U589  ( .A(\U1/aes_core/SB2/n2776 ), .Y(
        \U1/aes_core/SB2/n2874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U588  ( .A(\U1/aes_core/SB2/n2941 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2733 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U587  ( .A(\U1/aes_core/SB2/n2604 ), .Y(
        \U1/aes_core/SB2/n2910 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U586  ( .A(Dout[57]), .B(Dout[56]), .Y(
        \U1/aes_core/SB2/n2536 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U585  ( .A(\U1/aes_core/SB2/n2536 ), .B(
        \U1/aes_core/SB2/n2552 ), .Y(\U1/aes_core/SB2/n2842 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U584  ( .A(\U1/aes_core/SB2/n2842 ), .Y(
        \U1/aes_core/SB2/n2951 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U583  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2951 ), .Y(\U1/aes_core/SB2/n2847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U582  ( .A(\U1/aes_core/SB2/n2522 ), .B(
        Dout[57]), .Y(\U1/aes_core/SB2/n2551 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U581  ( .A(\U1/aes_core/SB2/n2533 ), .B(
        \U1/aes_core/SB2/n2551 ), .Y(\U1/aes_core/SB2/n2742 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U580  ( .A(\U1/aes_core/SB2/n2742 ), .Y(
        \U1/aes_core/SB2/n2831 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U579  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2711 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U578  ( .A(\U1/aes_core/SB2/n2733 ), .B(
        \U1/aes_core/SB2/n2847 ), .C(\U1/aes_core/SB2/n2711 ), .Y(
        \U1/aes_core/SB2/n2571 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U577  ( .A(\U1/aes_core/SB2/n2531 ), .B(
        \U1/aes_core/SB2/n2549 ), .Y(\U1/aes_core/SB2/n2775 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U576  ( .A(\U1/aes_core/SB2/n2523 ), .B(
        Dout[58]), .Y(\U1/aes_core/SB2/n2542 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U575  ( .A(\U1/aes_core/SB2/n2542 ), .B(
        \U1/aes_core/SB2/n2551 ), .Y(\U1/aes_core/SB2/n2773 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U574  ( .A(\U1/aes_core/SB2/n2775 ), .B(
        \U1/aes_core/SB2/n2773 ), .Y(\U1/aes_core/SB2/n2688 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U573  ( .A(\U1/aes_core/SB2/n2603 ), .Y(
        \U1/aes_core/SB2/n2912 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U572  ( .A(Dout[61]), .Y(
        \U1/aes_core/SB2/n2526 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U571  ( .A(\U1/aes_core/SB2/n2524 ), .B(
        \U1/aes_core/SB2/n2526 ), .Y(\U1/aes_core/SB2/n2550 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U570  ( .A(\U1/aes_core/SB2/n2540 ), .B(
        \U1/aes_core/SB2/n2550 ), .Y(\U1/aes_core/SB2/n2955 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U569  ( .A(\U1/aes_core/SB2/n2955 ), .Y(
        \U1/aes_core/SB2/n2865 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U568  ( .A(\U1/aes_core/SB2/n2525 ), .B(
        Dout[56]), .Y(\U1/aes_core/SB2/n2541 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U567  ( .A(\U1/aes_core/SB2/n2541 ), .B(
        \U1/aes_core/SB2/n2552 ), .Y(\U1/aes_core/SB2/n2920 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U566  ( .A(\U1/aes_core/SB2/n2920 ), .Y(
        \U1/aes_core/SB2/n2747 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U565  ( .A0(\U1/aes_core/SB2/n2912 ), 
        .A1(\U1/aes_core/SB2/n2865 ), .B0(\U1/aes_core/SB2/n2747 ), .Y(
        \U1/aes_core/SB2/n2530 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U564  ( .A(\U1/aes_core/SB2/n2536 ), .B(
        \U1/aes_core/SB2/n2533 ), .Y(\U1/aes_core/SB2/n2908 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U563  ( .A(\U1/aes_core/SB2/n2908 ), .Y(
        \U1/aes_core/SB2/n2873 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U562  ( .A(\U1/aes_core/SB2/n2526 ), .B(
        Dout[60]), .Y(\U1/aes_core/SB2/n2557 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U561  ( .A(\U1/aes_core/SB2/n2549 ), .B(
        \U1/aes_core/SB2/n2557 ), .Y(\U1/aes_core/SB2/n2948 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U560  ( .A(\U1/aes_core/SB2/n2775 ), .B(
        \U1/aes_core/SB2/n2948 ), .Y(\U1/aes_core/SB2/n2666 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U559  ( .A(\U1/aes_core/SB2/n2528 ), .B(
        \U1/aes_core/SB2/n2527 ), .Y(\U1/aes_core/SB2/n2548 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U558  ( .A(\U1/aes_core/SB2/n2539 ), .B(
        \U1/aes_core/SB2/n2548 ), .Y(\U1/aes_core/SB2/n2923 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U557  ( .A(\U1/aes_core/SB2/n2923 ), .Y(
        \U1/aes_core/SB2/n2647 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U556  ( .A0(\U1/aes_core/SB2/n2873 ), 
        .A1(\U1/aes_core/SB2/n2666 ), .B0(\U1/aes_core/SB2/n2647 ), .B1(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2529 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U555  ( .AN(\U1/aes_core/SB2/n2688 ), 
        .B(\U1/aes_core/SB2/n2530 ), .C(\U1/aes_core/SB2/n2529 ), .Y(
        \U1/aes_core/SB2/n2570 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U554  ( .A(\U1/aes_core/SB2/n2531 ), .B(
        \U1/aes_core/SB2/n2548 ), .Y(\U1/aes_core/SB2/n2792 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U553  ( .A(\U1/aes_core/SB2/n2535 ), .B(
        \U1/aes_core/SB2/n2536 ), .Y(\U1/aes_core/SB2/n2958 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U552  ( .A(\U1/aes_core/SB2/n2558 ), .B(
        \U1/aes_core/SB2/n2539 ), .Y(\U1/aes_core/SB2/n2843 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U551  ( .A(\U1/aes_core/SB2/n2535 ), .B(
        \U1/aes_core/SB2/n2541 ), .Y(\U1/aes_core/SB2/n2840 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U550  ( .A(\U1/aes_core/SB2/n2532 ), .B(
        \U1/aes_core/SB2/n2542 ), .Y(\U1/aes_core/SB2/n2845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U549  ( .A(\U1/aes_core/SB2/n2845 ), .Y(
        \U1/aes_core/SB2/n2825 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U548  ( .A(\U1/aes_core/SB2/n2948 ), .Y(
        \U1/aes_core/SB2/n2661 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U547  ( .A(\U1/aes_core/SB2/n2533 ), .B(
        \U1/aes_core/SB2/n2541 ), .Y(\U1/aes_core/SB2/n2863 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U546  ( .A(\U1/aes_core/SB2/n2863 ), .Y(
        \U1/aes_core/SB2/n2909 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U545  ( .A0(\U1/aes_core/SB2/n2825 ), 
        .A1(\U1/aes_core/SB2/n2910 ), .B0(\U1/aes_core/SB2/n2661 ), .B1(
        \U1/aes_core/SB2/n2909 ), .Y(\U1/aes_core/SB2/n2534 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U544  ( .A0(\U1/aes_core/SB2/n2792 ), 
        .A1(\U1/aes_core/SB2/n2958 ), .B0(\U1/aes_core/SB2/n2843 ), .B1(
        \U1/aes_core/SB2/n2840 ), .C0(\U1/aes_core/SB2/n2534 ), .Y(
        \U1/aes_core/SB2/n2569 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U543  ( .A(\U1/aes_core/SB2/n2845 ), .B(
        \U1/aes_core/SB2/n2792 ), .Y(\U1/aes_core/SB2/n2654 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U542  ( .A(\U1/aes_core/SB2/n2840 ), .B(
        \U1/aes_core/SB2/n2775 ), .Y(\U1/aes_core/SB2/n2664 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U541  ( .A(\U1/aes_core/SB2/n2664 ), .Y(
        \U1/aes_core/SB2/n2538 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U540  ( .A(\U1/aes_core/SB2/n2535 ), .B(
        \U1/aes_core/SB2/n2551 ), .Y(\U1/aes_core/SB2/n2936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U539  ( .A(\U1/aes_core/SB2/n2936 ), .Y(
        \U1/aes_core/SB2/n2864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U538  ( .A(\U1/aes_core/SB2/n2536 ), .B(
        \U1/aes_core/SB2/n2542 ), .Y(\U1/aes_core/SB2/n2921 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U537  ( .A(\U1/aes_core/SB2/n2921 ), .Y(
        \U1/aes_core/SB2/n2932 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U536  ( .A0(\U1/aes_core/SB2/n2864 ), 
        .A1(\U1/aes_core/SB2/n2932 ), .B0(\U1/aes_core/SB2/n2865 ), .Y(
        \U1/aes_core/SB2/n2537 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U535  ( .A(\U1/aes_core/SB2/n2540 ), .B(
        \U1/aes_core/SB2/n2557 ), .Y(\U1/aes_core/SB2/n2937 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U534  ( .A(\U1/aes_core/SB2/n2937 ), .Y(
        \U1/aes_core/SB2/n2866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U533  ( .A(\U1/aes_core/SB2/n2866 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2681 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U532  ( .AN(\U1/aes_core/SB2/n2654 ), 
        .B(\U1/aes_core/SB2/n2538 ), .C(\U1/aes_core/SB2/n2537 ), .D(
        \U1/aes_core/SB2/n2681 ), .Y(\U1/aes_core/SB2/n2547 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U531  ( .A(\U1/aes_core/SB2/n2550 ), .B(
        \U1/aes_core/SB2/n2548 ), .Y(\U1/aes_core/SB2/n2957 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U530  ( .A(\U1/aes_core/SB2/n2540 ), .B(
        \U1/aes_core/SB2/n2539 ), .Y(\U1/aes_core/SB2/n2949 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U529  ( .A0(\U1/aes_core/SB2/n2603 ), 
        .A1(\U1/aes_core/SB2/n2755 ), .B0(\U1/aes_core/SB2/n2957 ), .B1(
        \U1/aes_core/SB2/n2845 ), .C0(\U1/aes_core/SB2/n2949 ), .C1(
        \U1/aes_core/SB2/n2863 ), .Y(\U1/aes_core/SB2/n2546 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U528  ( .A(\U1/aes_core/SB2/n2908 ), .B(
        \U1/aes_core/SB2/n2603 ), .Y(\U1/aes_core/SB2/n2739 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U527  ( .A(\U1/aes_core/SB2/n2661 ), .B(
        \U1/aes_core/SB2/n2825 ), .Y(\U1/aes_core/SB2/n2692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U526  ( .A(\U1/aes_core/SB2/n2909 ), .B(
        \U1/aes_core/SB2/n2910 ), .Y(\U1/aes_core/SB2/n2712 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U525  ( .A(\U1/aes_core/SB2/n2843 ), .Y(
        \U1/aes_core/SB2/n2938 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U524  ( .A(\U1/aes_core/SB2/n2938 ), .B(
        \U1/aes_core/SB2/n2747 ), .Y(\U1/aes_core/SB2/n2750 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U523  ( .AN(\U1/aes_core/SB2/n2739 ), 
        .B(\U1/aes_core/SB2/n2692 ), .C(\U1/aes_core/SB2/n2712 ), .D(
        \U1/aes_core/SB2/n2750 ), .Y(\U1/aes_core/SB2/n2545 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U522  ( .A(\U1/aes_core/SB2/n2558 ), .B(
        \U1/aes_core/SB2/n2550 ), .Y(\U1/aes_core/SB2/n2662 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U521  ( .A(\U1/aes_core/SB2/n2662 ), .B(
        \U1/aes_core/SB2/n2920 ), .Y(\U1/aes_core/SB2/n2816 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U520  ( .A(\U1/aes_core/SB2/n2542 ), .B(
        \U1/aes_core/SB2/n2541 ), .Y(\U1/aes_core/SB2/n2956 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U519  ( .A(\U1/aes_core/SB2/n2923 ), .B(
        \U1/aes_core/SB2/n2956 ), .Y(\U1/aes_core/SB2/n2781 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U518  ( .A(\U1/aes_core/SB2/n2781 ), .Y(
        \U1/aes_core/SB2/n2543 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U517  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2747 ), .Y(\U1/aes_core/SB2/n2800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U516  ( .A(\U1/aes_core/SB2/n2956 ), .Y(
        \U1/aes_core/SB2/n2939 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U515  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2939 ), .Y(\U1/aes_core/SB2/n2851 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U514  ( .AN(\U1/aes_core/SB2/n2816 ), 
        .B(\U1/aes_core/SB2/n2543 ), .C(\U1/aes_core/SB2/n2800 ), .D(
        \U1/aes_core/SB2/n2851 ), .Y(\U1/aes_core/SB2/n2544 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U513  ( .A(\U1/aes_core/SB2/n2547 ), .B(
        \U1/aes_core/SB2/n2546 ), .C(\U1/aes_core/SB2/n2545 ), .D(
        \U1/aes_core/SB2/n2544 ), .Y(\U1/aes_core/SB2/n2643 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U512  ( .A(\U1/aes_core/SB2/n2842 ), .B(
        \U1/aes_core/SB2/n2662 ), .Y(\U1/aes_core/SB2/n2850 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U511  ( .A(\U1/aes_core/SB2/n2557 ), .B(
        \U1/aes_core/SB2/n2548 ), .Y(\U1/aes_core/SB2/n2758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U510  ( .A(\U1/aes_core/SB2/n2824 ), .B(
        \U1/aes_core/SB2/n2758 ), .Y(\U1/aes_core/SB2/n2729 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U509  ( .A(\U1/aes_core/SB2/n2957 ), .Y(
        \U1/aes_core/SB2/n2913 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U508  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2873 ), .Y(\U1/aes_core/SB2/n2678 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U507  ( .A0(\U1/aes_core/SB2/n2758 ), 
        .A1(\U1/aes_core/SB2/n2956 ), .B0(\U1/aes_core/SB2/n2678 ), .Y(
        \U1/aes_core/SB2/n2556 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U506  ( .A(\U1/aes_core/SB2/n2773 ), .Y(
        \U1/aes_core/SB2/n2868 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U505  ( .A(\U1/aes_core/SB2/n2868 ), .B(
        \U1/aes_core/SB2/n2912 ), .Y(\U1/aes_core/SB2/n2869 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U504  ( .A(\U1/aes_core/SB2/n2912 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2828 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U503  ( .A(\U1/aes_core/SB2/n2550 ), .B(
        \U1/aes_core/SB2/n2549 ), .Y(\U1/aes_core/SB2/n2919 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U502  ( .A(\U1/aes_core/SB2/n2919 ), .Y(
        \U1/aes_core/SB2/n2673 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U501  ( .A(\U1/aes_core/SB2/n2864 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2697 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U500  ( .A(\U1/aes_core/SB2/n2907 ), .Y(
        \U1/aes_core/SB2/n2867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U499  ( .A(\U1/aes_core/SB2/n2867 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2761 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U498  ( .A(\U1/aes_core/SB2/n2869 ), .B(
        \U1/aes_core/SB2/n2828 ), .C(\U1/aes_core/SB2/n2697 ), .D(
        \U1/aes_core/SB2/n2761 ), .Y(\U1/aes_core/SB2/n2555 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U497  ( .A(\U1/aes_core/SB2/n2909 ), .B(
        \U1/aes_core/SB2/n2866 ), .Y(\U1/aes_core/SB2/n2795 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U496  ( .A(\U1/aes_core/SB2/n2951 ), .B(
        \U1/aes_core/SB2/n2866 ), .Y(\U1/aes_core/SB2/n2786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U495  ( .A(\U1/aes_core/SB2/n2949 ), .Y(
        \U1/aes_core/SB2/n2942 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U494  ( .A(\U1/aes_core/SB2/n2825 ), .B(
        \U1/aes_core/SB2/n2942 ), .Y(\U1/aes_core/SB2/n2658 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U493  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2864 ), .Y(\U1/aes_core/SB2/n2769 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U492  ( .A(\U1/aes_core/SB2/n2795 ), .B(
        \U1/aes_core/SB2/n2786 ), .C(\U1/aes_core/SB2/n2658 ), .D(
        \U1/aes_core/SB2/n2769 ), .Y(\U1/aes_core/SB2/n2554 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U491  ( .A(\U1/aes_core/SB2/n2840 ), .Y(
        \U1/aes_core/SB2/n2809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U490  ( .A(\U1/aes_core/SB2/n2661 ), .B(
        \U1/aes_core/SB2/n2809 ), .Y(\U1/aes_core/SB2/n2645 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U489  ( .A(\U1/aes_core/SB2/n2552 ), .B(
        \U1/aes_core/SB2/n2551 ), .Y(\U1/aes_core/SB2/n2875 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U488  ( .A(\U1/aes_core/SB2/n2875 ), .Y(
        \U1/aes_core/SB2/n2930 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U487  ( .A(\U1/aes_core/SB2/n2661 ), .B(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2709 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U486  ( .A(\U1/aes_core/SB2/n2824 ), .Y(
        \U1/aes_core/SB2/n2953 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U485  ( .A(\U1/aes_core/SB2/n2953 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2744 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U484  ( .A(\U1/aes_core/SB2/n2865 ), .B(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2914 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U483  ( .A(\U1/aes_core/SB2/n2645 ), .B(
        \U1/aes_core/SB2/n2709 ), .C(\U1/aes_core/SB2/n2744 ), .D(
        \U1/aes_core/SB2/n2914 ), .Y(\U1/aes_core/SB2/n2553 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U482  ( .A(\U1/aes_core/SB2/n2850 ), .B(
        \U1/aes_core/SB2/n2729 ), .C(\U1/aes_core/SB2/n2556 ), .D(
        \U1/aes_core/SB2/n2555 ), .E(\U1/aes_core/SB2/n2554 ), .F(
        \U1/aes_core/SB2/n2553 ), .Y(\U1/aes_core/SB2/n2632 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U481  ( .A(\U1/aes_core/SB2/n2632 ), .Y(
        \U1/aes_core/SB2/n2567 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U480  ( .A(\U1/aes_core/SB2/n2921 ), .B(
        \U1/aes_core/SB2/n2758 ), .Y(\U1/aes_core/SB2/n2655 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U479  ( .A(\U1/aes_core/SB2/n2558 ), .B(
        \U1/aes_core/SB2/n2557 ), .Y(\U1/aes_core/SB2/n2918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U478  ( .A(\U1/aes_core/SB2/n2918 ), .B(
        \U1/aes_core/SB2/n2773 ), .Y(\U1/aes_core/SB2/n2782 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U477  ( .A(\U1/aes_core/SB2/n2782 ), .Y(
        \U1/aes_core/SB2/n2560 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U476  ( .A(\U1/aes_core/SB2/n2775 ), .Y(
        \U1/aes_core/SB2/n2943 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U475  ( .A0(\U1/aes_core/SB2/n2673 ), 
        .A1(\U1/aes_core/SB2/n2943 ), .B0(\U1/aes_core/SB2/n2930 ), .Y(
        \U1/aes_core/SB2/n2559 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U474  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2809 ), .Y(\U1/aes_core/SB2/n2680 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U473  ( .AN(\U1/aes_core/SB2/n2655 ), 
        .B(\U1/aes_core/SB2/n2560 ), .C(\U1/aes_core/SB2/n2559 ), .D(
        \U1/aes_core/SB2/n2680 ), .Y(\U1/aes_core/SB2/n2564 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U472  ( .A0(\U1/aes_core/SB2/n2907 ), 
        .A1(\U1/aes_core/SB2/n2955 ), .B0(\U1/aes_core/SB2/n2792 ), .B1(
        \U1/aes_core/SB2/n2840 ), .C0(\U1/aes_core/SB2/n2920 ), .C1(
        \U1/aes_core/SB2/n2937 ), .Y(\U1/aes_core/SB2/n2563 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U471  ( .A(\U1/aes_core/SB2/n2955 ), .B(
        \U1/aes_core/SB2/n2958 ), .Y(\U1/aes_core/SB2/n2720 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U470  ( .A(\U1/aes_core/SB2/n2943 ), .B(
        \U1/aes_core/SB2/n2864 ), .Y(\U1/aes_core/SB2/n2853 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U469  ( .A(\U1/aes_core/SB2/n2825 ), .B(
        \U1/aes_core/SB2/n2943 ), .Y(\U1/aes_core/SB2/n2787 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U468  ( .A(\U1/aes_core/SB2/n2809 ), .B(
        \U1/aes_core/SB2/n2910 ), .Y(\U1/aes_core/SB2/n2659 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U467  ( .AN(\U1/aes_core/SB2/n2720 ), 
        .B(\U1/aes_core/SB2/n2853 ), .C(\U1/aes_core/SB2/n2787 ), .D(
        \U1/aes_core/SB2/n2659 ), .Y(\U1/aes_core/SB2/n2562 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U466  ( .A(\U1/aes_core/SB2/n2953 ), .B(
        \U1/aes_core/SB2/n2938 ), .Y(\U1/aes_core/SB2/n2732 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U465  ( .A(\U1/aes_core/SB2/n2809 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U464  ( .A(\U1/aes_core/SB2/n2661 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U463  ( .A(\U1/aes_core/SB2/n2868 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2745 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U462  ( .A(\U1/aes_core/SB2/n2732 ), .B(
        \U1/aes_core/SB2/n2799 ), .C(\U1/aes_core/SB2/n2700 ), .D(
        \U1/aes_core/SB2/n2745 ), .Y(\U1/aes_core/SB2/n2561 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U461  ( .A(\U1/aes_core/SB2/n2564 ), .B(
        \U1/aes_core/SB2/n2563 ), .C(\U1/aes_core/SB2/n2562 ), .D(
        \U1/aes_core/SB2/n2561 ), .Y(\U1/aes_core/SB2/n2565 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U460  ( .A(\U1/aes_core/SB2/n2565 ), .Y(
        \U1/aes_core/SB2/n2935 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U459  ( .A(\U1/aes_core/SB2/n2951 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2566 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U458  ( .AN(\U1/aes_core/SB2/n2643 ), 
        .B(\U1/aes_core/SB2/n2567 ), .C(\U1/aes_core/SB2/n2935 ), .D(
        \U1/aes_core/SB2/n2566 ), .Y(\U1/aes_core/SB2/n2568 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U457  ( .A(\U1/aes_core/SB2/n2693 ), .B(
        \U1/aes_core/SB2/n2790 ), .C(\U1/aes_core/SB2/n2571 ), .D(
        \U1/aes_core/SB2/n2570 ), .E(\U1/aes_core/SB2/n2569 ), .F(
        \U1/aes_core/SB2/n2568 ), .Y(\U1/aes_core/SB2/n2622 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U456  ( .A(\U1/aes_core/SB2/n2936 ), .B(
        \U1/aes_core/SB2/n2603 ), .Y(\U1/aes_core/SB2/n2738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U455  ( .A(\U1/aes_core/SB2/n2865 ), .B(
        \U1/aes_core/SB2/n2953 ), .Y(\U1/aes_core/SB2/n2789 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U454  ( .A(\U1/aes_core/SB2/n2942 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2691 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U453  ( .A(\U1/aes_core/SB2/n2662 ), .Y(
        \U1/aes_core/SB2/n2931 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U452  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2714 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U451  ( .AN(\U1/aes_core/SB2/n2738 ), 
        .B(\U1/aes_core/SB2/n2789 ), .C(\U1/aes_core/SB2/n2691 ), .D(
        \U1/aes_core/SB2/n2714 ), .Y(\U1/aes_core/SB2/n2578 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U450  ( .A(\U1/aes_core/SB2/n2923 ), .B(
        \U1/aes_core/SB2/n2773 ), .Y(\U1/aes_core/SB2/n2815 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U449  ( .A(\U1/aes_core/SB2/n2825 ), .B(
        \U1/aes_core/SB2/n2912 ), .Y(\U1/aes_core/SB2/n2671 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U448  ( .A0(\U1/aes_core/SB2/n2932 ), 
        .A1(\U1/aes_core/SB2/n2831 ), .B0(\U1/aes_core/SB2/n2661 ), .Y(
        \U1/aes_core/SB2/n2572 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U447  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2763 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U446  ( .AN(\U1/aes_core/SB2/n2815 ), 
        .B(\U1/aes_core/SB2/n2671 ), .C(\U1/aes_core/SB2/n2572 ), .D(
        \U1/aes_core/SB2/n2763 ), .Y(\U1/aes_core/SB2/n2573 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U445  ( .A(\U1/aes_core/SB2/n2573 ), .Y(
        \U1/aes_core/SB2/n2577 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U444  ( .A(\U1/aes_core/SB2/n2792 ), .Y(
        \U1/aes_core/SB2/n2933 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U443  ( .A(\U1/aes_core/SB2/n2958 ), .Y(
        \U1/aes_core/SB2/n2832 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U442  ( .A0(\U1/aes_core/SB2/n2953 ), 
        .A1(\U1/aes_core/SB2/n2866 ), .B0(\U1/aes_core/SB2/n2933 ), .B1(
        \U1/aes_core/SB2/n2747 ), .C0(\U1/aes_core/SB2/n2832 ), .C1(
        \U1/aes_core/SB2/n2931 ), .Y(\U1/aes_core/SB2/n2576 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U441  ( .A0(\U1/aes_core/SB2/n2758 ), 
        .A1(\U1/aes_core/SB2/n2936 ), .B0(\U1/aes_core/SB2/n2956 ), .B1(
        \U1/aes_core/SB2/n2957 ), .Y(\U1/aes_core/SB2/n2574 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U440  ( .A0(\U1/aes_core/SB2/n2809 ), 
        .A1(\U1/aes_core/SB2/n2647 ), .B0(\U1/aes_core/SB2/n2865 ), .B1(
        \U1/aes_core/SB2/n2909 ), .C0(\U1/aes_core/SB2/n2574 ), .Y(
        \U1/aes_core/SB2/n2575 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U439  ( .AN(\U1/aes_core/SB2/n2578 ), 
        .B(\U1/aes_core/SB2/n2577 ), .C(\U1/aes_core/SB2/n2576 ), .D(
        \U1/aes_core/SB2/n2575 ), .Y(\U1/aes_core/SB2/n2641 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U438  ( .A(\U1/aes_core/SB2/n2957 ), .B(
        \U1/aes_core/SB2/n2773 ), .Y(\U1/aes_core/SB2/n2656 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U437  ( .A0(\U1/aes_core/SB2/n2843 ), 
        .A1(\U1/aes_core/SB2/n2957 ), .B0(\U1/aes_core/SB2/n2875 ), .Y(
        \U1/aes_core/SB2/n2583 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U436  ( .A(\U1/aes_core/SB2/n2875 ), .B(
        \U1/aes_core/SB2/n2863 ), .Y(\U1/aes_core/SB2/n2740 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB2/U435  ( .A0(\U1/aes_core/SB2/n2864 ), .A1(
        \U1/aes_core/SB2/n2647 ), .B0(\U1/aes_core/SB2/n2740 ), .B1(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2582 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U434  ( .A0(\U1/aes_core/SB2/n2918 ), 
        .A1(\U1/aes_core/SB2/n2958 ), .B0(\U1/aes_core/SB2/n2662 ), .B1(
        \U1/aes_core/SB2/n2755 ), .C0(\U1/aes_core/SB2/n2920 ), .C1(
        \U1/aes_core/SB2/n2949 ), .Y(\U1/aes_core/SB2/n2581 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U433  ( .A(\U1/aes_core/SB2/n2758 ), .Y(
        \U1/aes_core/SB2/n2826 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U432  ( .A(\U1/aes_core/SB2/n2951 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2852 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U431  ( .A(\U1/aes_core/SB2/n2825 ), .B(
        \U1/aes_core/SB2/n2647 ), .Y(\U1/aes_core/SB2/n2679 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U430  ( .A(\U1/aes_core/SB2/n2661 ), .B(
        \U1/aes_core/SB2/n2868 ), .Y(\U1/aes_core/SB2/n2699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U429  ( .A(\U1/aes_core/SB2/n2825 ), .B(
        \U1/aes_core/SB2/n2866 ), .Y(\U1/aes_core/SB2/n2798 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U428  ( .A(\U1/aes_core/SB2/n2852 ), .B(
        \U1/aes_core/SB2/n2679 ), .C(\U1/aes_core/SB2/n2699 ), .D(
        \U1/aes_core/SB2/n2798 ), .Y(\U1/aes_core/SB2/n2580 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U427  ( .A(\U1/aes_core/SB2/n2845 ), .B(
        \U1/aes_core/SB2/n2758 ), .Y(\U1/aes_core/SB2/n2721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U426  ( .A(\U1/aes_core/SB2/n2831 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2731 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U425  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2747 ), .Y(\U1/aes_core/SB2/n2762 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB2/U424  ( .AN(\U1/aes_core/SB2/n2721 ), 
        .B(\U1/aes_core/SB2/n2731 ), .C(\U1/aes_core/SB2/n2762 ), .Y(
        \U1/aes_core/SB2/n2579 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U423  ( .A(\U1/aes_core/SB2/n2656 ), .B(
        \U1/aes_core/SB2/n2583 ), .C(\U1/aes_core/SB2/n2582 ), .D(
        \U1/aes_core/SB2/n2581 ), .E(\U1/aes_core/SB2/n2580 ), .F(
        \U1/aes_core/SB2/n2579 ), .Y(\U1/aes_core/SB2/n2964 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U422  ( .A0(\U1/aes_core/SB2/n2661 ), 
        .A1(\U1/aes_core/SB2/n2910 ), .B0(\U1/aes_core/SB2/n2941 ), .Y(
        \U1/aes_core/SB2/n2584 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U421  ( .A(\U1/aes_core/SB2/n2647 ), .B(
        \U1/aes_core/SB2/n2747 ), .Y(\U1/aes_core/SB2/n2784 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U420  ( .A(\U1/aes_core/SB2/n2864 ), .B(
        \U1/aes_core/SB2/n2933 ), .Y(\U1/aes_core/SB2/n2676 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U419  ( .A(\U1/aes_core/SB2/n2933 ), .B(
        \U1/aes_core/SB2/n2868 ), .Y(\U1/aes_core/SB2/n2727 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U418  ( .A(\U1/aes_core/SB2/n2584 ), .B(
        \U1/aes_core/SB2/n2784 ), .C(\U1/aes_core/SB2/n2676 ), .D(
        \U1/aes_core/SB2/n2727 ), .Y(\U1/aes_core/SB2/n2588 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U417  ( .A0(\U1/aes_core/SB2/n2936 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2662 ), .B1(
        \U1/aes_core/SB2/n2908 ), .C0(\U1/aes_core/SB2/n2937 ), .C1(
        \U1/aes_core/SB2/n2773 ), .Y(\U1/aes_core/SB2/n2587 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U416  ( .A(\U1/aes_core/SB2/n2867 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U415  ( .A(\U1/aes_core/SB2/n2866 ), .B(
        \U1/aes_core/SB2/n2939 ), .Y(\U1/aes_core/SB2/n2848 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U414  ( .A(\U1/aes_core/SB2/n2866 ), .B(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2695 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U413  ( .A(\U1/aes_core/SB2/n2942 ), .B(
        \U1/aes_core/SB2/n2932 ), .Y(\U1/aes_core/SB2/n2657 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U412  ( .A(\U1/aes_core/SB2/n2708 ), .B(
        \U1/aes_core/SB2/n2848 ), .C(\U1/aes_core/SB2/n2695 ), .D(
        \U1/aes_core/SB2/n2657 ), .Y(\U1/aes_core/SB2/n2586 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U411  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2770 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U410  ( .A(\U1/aes_core/SB2/n2951 ), .B(
        \U1/aes_core/SB2/n2912 ), .Y(\U1/aes_core/SB2/n2743 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U409  ( .A(\U1/aes_core/SB2/n2941 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2794 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U408  ( .A(\U1/aes_core/SB2/n2673 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2644 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U407  ( .A(\U1/aes_core/SB2/n2770 ), .B(
        \U1/aes_core/SB2/n2743 ), .C(\U1/aes_core/SB2/n2794 ), .D(
        \U1/aes_core/SB2/n2644 ), .Y(\U1/aes_core/SB2/n2585 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U406  ( .A(\U1/aes_core/SB2/n2588 ), .B(
        \U1/aes_core/SB2/n2587 ), .C(\U1/aes_core/SB2/n2586 ), .D(
        \U1/aes_core/SB2/n2585 ), .Y(\U1/aes_core/SB2/n2630 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U405  ( .A(\U1/aes_core/SB2/n2622 ), .B(
        \U1/aes_core/SB2/n2641 ), .C(\U1/aes_core/SB2/n2964 ), .D(
        \U1/aes_core/SB2/n2630 ), .Y(\U1/aes_core/SB2/n2597 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U404  ( .A(\U1/aes_core/SB2/n2918 ), .Y(
        \U1/aes_core/SB2/n2821 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U403  ( .A0(\U1/aes_core/SB2/n2773 ), 
        .A1(\U1/aes_core/SB2/n2604 ), .B0(\U1/aes_core/SB2/n2742 ), .B1(
        \U1/aes_core/SB2/n2949 ), .Y(\U1/aes_core/SB2/n2589 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U402  ( .A0(\U1/aes_core/SB2/n2821 ), 
        .A1(\U1/aes_core/SB2/n2873 ), .B0(\U1/aes_core/SB2/n2943 ), .B1(
        \U1/aes_core/SB2/n2951 ), .C0(\U1/aes_core/SB2/n2589 ), .Y(
        \U1/aes_core/SB2/n2596 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U401  ( .A(\U1/aes_core/SB2/n2842 ), .B(
        \U1/aes_core/SB2/n2845 ), .Y(\U1/aes_core/SB2/n2841 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U400  ( .A0(\U1/aes_core/SB2/n2776 ), 
        .A1(\U1/aes_core/SB2/n2845 ), .B0(\U1/aes_core/SB2/n2758 ), .B1(
        \U1/aes_core/SB2/n2907 ), .Y(\U1/aes_core/SB2/n2590 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U399  ( .A0(\U1/aes_core/SB2/n2673 ), 
        .A1(\U1/aes_core/SB2/n2841 ), .B0(\U1/aes_core/SB2/n2913 ), .B1(
        \U1/aes_core/SB2/n2932 ), .C0(\U1/aes_core/SB2/n2590 ), .Y(
        \U1/aes_core/SB2/n2595 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U398  ( .A(\U1/aes_core/SB2/n2937 ), .B(
        \U1/aes_core/SB2/n2775 ), .Y(\U1/aes_core/SB2/n2593 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U397  ( .A(\U1/aes_core/SB2/n2866 ), .B(
        \U1/aes_core/SB2/n2912 ), .Y(\U1/aes_core/SB2/n2833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U396  ( .A(\U1/aes_core/SB2/n2833 ), .Y(
        \U1/aes_core/SB2/n2592 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U395  ( .A(\U1/aes_core/SB2/n2824 ), .B(
        \U1/aes_core/SB2/n2918 ), .Y(\U1/aes_core/SB2/n2705 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U394  ( .A(\U1/aes_core/SB2/n2923 ), .B(
        \U1/aes_core/SB2/n2921 ), .Y(\U1/aes_core/SB2/n2858 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U392  ( .A(\U1/aes_core/SB2/n2873 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2715 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U390  ( .A0(\U1/aes_core/SB2/n2832 ), 
        .A1(\U1/aes_core/SB2/n2593 ), .B0(\U1/aes_core/SB2/n2809 ), .B1(
        \U1/aes_core/SB2/n2592 ), .C0(\U1/aes_core/SB2/n2591 ), .Y(
        \U1/aes_core/SB2/n2594 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U389  ( .AN(\U1/aes_core/SB2/n2597 ), 
        .B(\U1/aes_core/SB2/n2596 ), .C(\U1/aes_core/SB2/n2595 ), .D(
        \U1/aes_core/SB2/n2594 ), .Y(\U1/aes_core/sb2 [24]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U388  ( .A(\U1/aes_core/SB2/n2845 ), .B(
        \U1/aes_core/SB2/n2662 ), .Y(\U1/aes_core/SB2/n2722 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U387  ( .A(\U1/aes_core/SB2/n2792 ), .B(
        \U1/aes_core/SB2/n2842 ), .Y(\U1/aes_core/SB2/n2682 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U386  ( .A(\U1/aes_core/SB2/n2809 ), .B(
        \U1/aes_core/SB2/n2941 ), .Y(\U1/aes_core/SB2/n2791 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U385  ( .A0(\U1/aes_core/SB2/n2791 ), 
        .A1(\U1/aes_core/SB2/n2845 ), .B0(\U1/aes_core/SB2/n2955 ), .Y(
        \U1/aes_core/SB2/n2602 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U384  ( .A(\U1/aes_core/SB2/n2873 ), .B(
        \U1/aes_core/SB2/n2942 ), .Y(\U1/aes_core/SB2/n2698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U383  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2873 ), .Y(\U1/aes_core/SB2/n2797 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U382  ( .A(\U1/aes_core/SB2/n2939 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2730 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U381  ( .A(\U1/aes_core/SB2/n2698 ), .B(
        \U1/aes_core/SB2/n2797 ), .C(\U1/aes_core/SB2/n2730 ), .Y(
        \U1/aes_core/SB2/n2601 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U380  ( .A(\U1/aes_core/SB2/n2873 ), .B(
        \U1/aes_core/SB2/n2953 ), .Y(\U1/aes_core/SB2/n2757 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U379  ( .A(\U1/aes_core/SB2/n2939 ), .B(
        \U1/aes_core/SB2/n2930 ), .C(\U1/aes_core/SB2/n2951 ), .Y(
        \U1/aes_core/SB2/n2598 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U378  ( .A0(\U1/aes_core/SB2/n2757 ), 
        .A1(\U1/aes_core/SB2/n2919 ), .B0(\U1/aes_core/SB2/n2598 ), .B1(
        \U1/aes_core/SB2/n2949 ), .C0(\U1/aes_core/SB2/n2792 ), .C1(
        \U1/aes_core/SB2/n2824 ), .Y(\U1/aes_core/SB2/n2600 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U377  ( .A0(\U1/aes_core/SB2/n2920 ), 
        .A1(\U1/aes_core/SB2/n2948 ), .B0(\U1/aes_core/SB2/n2921 ), .B1(
        \U1/aes_core/SB2/n2918 ), .Y(\U1/aes_core/SB2/n2599 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U376  ( .A(\U1/aes_core/SB2/n2722 ), .B(
        \U1/aes_core/SB2/n2682 ), .C(\U1/aes_core/SB2/n2602 ), .D(
        \U1/aes_core/SB2/n2601 ), .E(\U1/aes_core/SB2/n2600 ), .F(
        \U1/aes_core/SB2/n2599 ), .Y(\U1/aes_core/SB2/n2963 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U375  ( .A(\U1/aes_core/SB2/n2773 ), .B(
        \U1/aes_core/SB2/n2758 ), .Y(\U1/aes_core/SB2/n2648 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U374  ( .A0(\U1/aes_core/SB2/n2773 ), 
        .A1(\U1/aes_core/SB2/n2863 ), .B0(\U1/aes_core/SB2/n2662 ), .Y(
        \U1/aes_core/SB2/n2609 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U373  ( .A(\U1/aes_core/SB2/n2867 ), .B(
        \U1/aes_core/SB2/n2873 ), .Y(\U1/aes_core/SB2/n2650 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U372  ( .A0(\U1/aes_core/SB2/n2755 ), 
        .A1(\U1/aes_core/SB2/n2923 ), .B0(\U1/aes_core/SB2/n2650 ), .B1(
        \U1/aes_core/SB2/n2937 ), .Y(\U1/aes_core/SB2/n2608 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U371  ( .A0(\U1/aes_core/SB2/n2742 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2907 ), .B1(
        \U1/aes_core/SB2/n2792 ), .C0(\U1/aes_core/SB2/n2921 ), .C1(
        \U1/aes_core/SB2/n2843 ), .Y(\U1/aes_core/SB2/n2607 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U370  ( .A(\U1/aes_core/SB2/n2956 ), .B(
        \U1/aes_core/SB2/n2603 ), .Y(\U1/aes_core/SB2/n2706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U369  ( .A(\U1/aes_core/SB2/n2943 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U368  ( .A(\U1/aes_core/SB2/n2864 ), .B(
        \U1/aes_core/SB2/n2938 ), .Y(\U1/aes_core/SB2/n2723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U367  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2953 ), .Y(\U1/aes_core/SB2/n2827 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U366  ( .AN(\U1/aes_core/SB2/n2706 ), 
        .B(\U1/aes_core/SB2/n2713 ), .C(\U1/aes_core/SB2/n2723 ), .D(
        \U1/aes_core/SB2/n2827 ), .Y(\U1/aes_core/SB2/n2606 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U365  ( .A(\U1/aes_core/SB2/n2824 ), .B(
        \U1/aes_core/SB2/n2604 ), .Y(\U1/aes_core/SB2/n2806 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U364  ( .A(\U1/aes_core/SB2/n2923 ), .B(
        \U1/aes_core/SB2/n2907 ), .Y(\U1/aes_core/SB2/n2859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U362  ( .A(\U1/aes_core/SB2/n2647 ), .B(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2672 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U360  ( .A(\U1/aes_core/SB2/n2648 ), .B(
        \U1/aes_core/SB2/n2609 ), .C(\U1/aes_core/SB2/n2608 ), .D(
        \U1/aes_core/SB2/n2607 ), .E(\U1/aes_core/SB2/n2606 ), .F(
        \U1/aes_core/SB2/n2605 ), .Y(\U1/aes_core/SB2/n2642 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U359  ( .A(\U1/aes_core/SB2/n2840 ), .B(
        \U1/aes_core/SB2/n2662 ), .Y(\U1/aes_core/SB2/n2660 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U358  ( .A(\U1/aes_core/SB2/n2792 ), .B(
        \U1/aes_core/SB2/n2742 ), .Y(\U1/aes_core/SB2/n2872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U357  ( .A(\U1/aes_core/SB2/n2773 ), .B(
        \U1/aes_core/SB2/n2843 ), .Y(\U1/aes_core/SB2/n2710 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U356  ( .A(\U1/aes_core/SB2/n2958 ), .B(
        \U1/aes_core/SB2/n2843 ), .Y(\U1/aes_core/SB2/n2725 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U355  ( .A(\U1/aes_core/SB2/n2868 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2785 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U354  ( .A(\U1/aes_core/SB2/n2939 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2677 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U353  ( .A(\U1/aes_core/SB2/n2943 ), .B(
        \U1/aes_core/SB2/n2939 ), .Y(\U1/aes_core/SB2/n2771 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U352  ( .A(\U1/aes_core/SB2/n2832 ), .B(
        \U1/aes_core/SB2/n2910 ), .Y(\U1/aes_core/SB2/n2696 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U351  ( .A(\U1/aes_core/SB2/n2785 ), .B(
        \U1/aes_core/SB2/n2677 ), .C(\U1/aes_core/SB2/n2771 ), .D(
        \U1/aes_core/SB2/n2696 ), .Y(\U1/aes_core/SB2/n2613 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U350  ( .A(\U1/aes_core/SB2/n2958 ), .B(
        \U1/aes_core/SB2/n2758 ), .Y(\U1/aes_core/SB2/n2746 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U349  ( .A(\U1/aes_core/SB2/n2957 ), .B(
        \U1/aes_core/SB2/n2742 ), .Y(\U1/aes_core/SB2/n2846 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U348  ( .A(\U1/aes_core/SB2/n2863 ), .B(
        \U1/aes_core/SB2/n2923 ), .Y(\U1/aes_core/SB2/n2796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U347  ( .A(\U1/aes_core/SB2/n2824 ), .B(
        \U1/aes_core/SB2/n2923 ), .Y(\U1/aes_core/SB2/n2646 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U346  ( .A0(\U1/aes_core/SB2/n2923 ), 
        .A1(\U1/aes_core/SB2/n2958 ), .B0(\U1/aes_core/SB2/n2758 ), .B1(
        \U1/aes_core/SB2/n2863 ), .Y(\U1/aes_core/SB2/n2611 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U345  ( .A0(\U1/aes_core/SB2/n2742 ), 
        .A1(\U1/aes_core/SB2/n2955 ), .B0(\U1/aes_core/SB2/n2755 ), .B1(
        \U1/aes_core/SB2/n2792 ), .Y(\U1/aes_core/SB2/n2610 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U344  ( .A(\U1/aes_core/SB2/n2746 ), .B(
        \U1/aes_core/SB2/n2846 ), .C(\U1/aes_core/SB2/n2796 ), .D(
        \U1/aes_core/SB2/n2646 ), .E(\U1/aes_core/SB2/n2611 ), .F(
        \U1/aes_core/SB2/n2610 ), .Y(\U1/aes_core/SB2/n2612 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U343  ( .A(\U1/aes_core/SB2/n2660 ), .B(
        \U1/aes_core/SB2/n2872 ), .C(\U1/aes_core/SB2/n2710 ), .D(
        \U1/aes_core/SB2/n2725 ), .E(\U1/aes_core/SB2/n2613 ), .F(
        \U1/aes_core/SB2/n2612 ), .Y(\U1/aes_core/SB2/n2631 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U342  ( .A0(\U1/aes_core/SB2/n2868 ), 
        .A1(\U1/aes_core/SB2/n2865 ), .B0(\U1/aes_core/SB2/n2942 ), .B1(
        \U1/aes_core/SB2/n2809 ), .C0(\U1/aes_core/SB2/n2631 ), .Y(
        \U1/aes_core/SB2/n2614 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U341  ( .A(\U1/aes_core/SB2/n2614 ), .Y(
        \U1/aes_core/SB2/n2621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U340  ( .A(\U1/aes_core/SB2/n2921 ), .B(
        \U1/aes_core/SB2/n2863 ), .Y(\U1/aes_core/SB2/n2911 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U339  ( .A0(\U1/aes_core/SB2/n2867 ), 
        .A1(\U1/aes_core/SB2/n2911 ), .B0(\U1/aes_core/SB2/n2943 ), .Y(
        \U1/aes_core/SB2/n2617 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U338  ( .A0(\U1/aes_core/SB2/n2832 ), 
        .A1(\U1/aes_core/SB2/n2932 ), .B0(\U1/aes_core/SB2/n2874 ), .Y(
        \U1/aes_core/SB2/n2616 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U337  ( .A0(\U1/aes_core/SB2/n2831 ), 
        .A1(\U1/aes_core/SB2/n2873 ), .B0(\U1/aes_core/SB2/n2938 ), .Y(
        \U1/aes_core/SB2/n2615 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U336  ( .A(\U1/aes_core/SB2/n2864 ), .B(
        \U1/aes_core/SB2/n2931 ), .Y(\U1/aes_core/SB2/n2689 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U335  ( .A(\U1/aes_core/SB2/n2617 ), .B(
        \U1/aes_core/SB2/n2616 ), .C(\U1/aes_core/SB2/n2615 ), .D(
        \U1/aes_core/SB2/n2689 ), .Y(\U1/aes_core/SB2/n2620 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U334  ( .A(\U1/aes_core/SB2/n2930 ), .B(
        \U1/aes_core/SB2/n2825 ), .Y(\U1/aes_core/SB2/n2879 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB2/U333  ( .A(\U1/aes_core/SB2/n2879 ), .B(
        \U1/aes_core/SB2/n2920 ), .C(\U1/aes_core/SB2/n2907 ), .Y(
        \U1/aes_core/SB2/n2618 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U332  ( .A0(\U1/aes_core/SB2/n2863 ), 
        .A1(\U1/aes_core/SB2/n2957 ), .B0(\U1/aes_core/SB2/n2618 ), .B1(
        \U1/aes_core/SB2/n2918 ), .C0(\U1/aes_core/SB2/n2956 ), .C1(
        \U1/aes_core/SB2/n2948 ), .Y(\U1/aes_core/SB2/n2619 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U331  ( .A(\U1/aes_core/SB2/n2963 ), .B(
        \U1/aes_core/SB2/n2642 ), .C(\U1/aes_core/SB2/n2622 ), .D(
        \U1/aes_core/SB2/n2621 ), .E(\U1/aes_core/SB2/n2620 ), .F(
        \U1/aes_core/SB2/n2619 ), .Y(\U1/aes_core/sb2 [25]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U330  ( .A0(\U1/aes_core/SB2/n2912 ), 
        .A1(\U1/aes_core/SB2/n2932 ), .B0(\U1/aes_core/SB2/n2953 ), .B1(
        \U1/aes_core/SB2/n2943 ), .Y(\U1/aes_core/SB2/n2623 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U329  ( .A0(\U1/aes_core/SB2/n2842 ), 
        .A1(\U1/aes_core/SB2/n2957 ), .B0(\U1/aes_core/SB2/n2792 ), .B1(
        \U1/aes_core/SB2/n2863 ), .C0(\U1/aes_core/SB2/n2623 ), .Y(
        \U1/aes_core/SB2/n2629 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U328  ( .A(\U1/aes_core/SB2/n2938 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2726 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U327  ( .A(\U1/aes_core/SB2/n2912 ), .B(
        \U1/aes_core/SB2/n2867 ), .Y(\U1/aes_core/SB2/n2707 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U326  ( .A(\U1/aes_core/SB2/n2932 ), .B(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2675 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U325  ( .A(\U1/aes_core/SB2/n2831 ), .B(
        \U1/aes_core/SB2/n2874 ), .Y(\U1/aes_core/SB2/n2694 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U324  ( .A(\U1/aes_core/SB2/n2726 ), .B(
        \U1/aes_core/SB2/n2707 ), .C(\U1/aes_core/SB2/n2675 ), .D(
        \U1/aes_core/SB2/n2694 ), .Y(\U1/aes_core/SB2/n2628 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U323  ( .A(\U1/aes_core/SB2/n2958 ), .B(
        \U1/aes_core/SB2/n2936 ), .Y(\U1/aes_core/SB2/n2820 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U322  ( .A0(\U1/aes_core/SB2/n2868 ), 
        .A1(\U1/aes_core/SB2/n2820 ), .B0(\U1/aes_core/SB2/n2942 ), .Y(
        \U1/aes_core/SB2/n2626 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U321  ( .A0(\U1/aes_core/SB2/n2939 ), 
        .A1(\U1/aes_core/SB2/n2809 ), .B0(\U1/aes_core/SB2/n2821 ), .Y(
        \U1/aes_core/SB2/n2625 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U320  ( .A0(\U1/aes_core/SB2/n2826 ), 
        .A1(\U1/aes_core/SB2/n2866 ), .B0(\U1/aes_core/SB2/n2941 ), .Y(
        \U1/aes_core/SB2/n2624 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U319  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2939 ), .Y(\U1/aes_core/SB2/n2793 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U318  ( .A(\U1/aes_core/SB2/n2626 ), .B(
        \U1/aes_core/SB2/n2625 ), .C(\U1/aes_core/SB2/n2624 ), .D(
        \U1/aes_core/SB2/n2793 ), .Y(\U1/aes_core/SB2/n2627 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U317  ( .A(\U1/aes_core/SB2/n2632 ), .B(
        \U1/aes_core/SB2/n2631 ), .C(\U1/aes_core/SB2/n2630 ), .D(
        \U1/aes_core/SB2/n2629 ), .E(\U1/aes_core/SB2/n2628 ), .F(
        \U1/aes_core/SB2/n2627 ), .Y(\U1/aes_core/SB2/n2962 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U316  ( .A0(\U1/aes_core/SB2/n2747 ), 
        .A1(\U1/aes_core/SB2/n2943 ), .B0(\U1/aes_core/SB2/n2951 ), .B1(
        \U1/aes_core/SB2/n2865 ), .C0(\U1/aes_core/SB2/n2962 ), .Y(
        \U1/aes_core/SB2/n2633 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U315  ( .A(\U1/aes_core/SB2/n2633 ), .Y(
        \U1/aes_core/SB2/n2640 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U314  ( .A(\U1/aes_core/SB2/n2874 ), .B(
        \U1/aes_core/SB2/n2661 ), .Y(\U1/aes_core/SB2/n2783 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U313  ( .A1N(\U1/aes_core/SB2/n2783 ), 
        .A0(\U1/aes_core/SB2/n2913 ), .B0(\U1/aes_core/SB2/n2864 ), .Y(
        \U1/aes_core/SB2/n2636 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U312  ( .A0(\U1/aes_core/SB2/n2832 ), 
        .A1(\U1/aes_core/SB2/n2740 ), .B0(\U1/aes_core/SB2/n2912 ), .Y(
        \U1/aes_core/SB2/n2635 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U311  ( .A0(\U1/aes_core/SB2/n2939 ), 
        .A1(\U1/aes_core/SB2/n2873 ), .B0(\U1/aes_core/SB2/n2933 ), .Y(
        \U1/aes_core/SB2/n2634 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U310  ( .A(\U1/aes_core/SB2/n2910 ), .B(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2690 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U309  ( .A(\U1/aes_core/SB2/n2636 ), .B(
        \U1/aes_core/SB2/n2635 ), .C(\U1/aes_core/SB2/n2634 ), .D(
        \U1/aes_core/SB2/n2690 ), .Y(\U1/aes_core/SB2/n2639 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U308  ( .A(\U1/aes_core/SB2/n2909 ), .B(
        \U1/aes_core/SB2/n2941 ), .Y(\U1/aes_core/SB2/n2940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U307  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2866 ), .Y(\U1/aes_core/SB2/n2637 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U306  ( .A0(\U1/aes_core/SB2/n2940 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2637 ), .B1(
        \U1/aes_core/SB2/n2921 ), .C0(\U1/aes_core/SB2/n2843 ), .C1(
        \U1/aes_core/SB2/n2845 ), .Y(\U1/aes_core/SB2/n2638 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U305  ( .A(\U1/aes_core/SB2/n2643 ), .B(
        \U1/aes_core/SB2/n2642 ), .C(\U1/aes_core/SB2/n2641 ), .D(
        \U1/aes_core/SB2/n2640 ), .E(\U1/aes_core/SB2/n2639 ), .F(
        \U1/aes_core/SB2/n2638 ), .Y(\U1/aes_core/sb2 [26]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U304  ( .A(\U1/aes_core/SB2/n2747 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2945 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U303  ( .AN(\U1/aes_core/SB2/n2646 ), 
        .B(\U1/aes_core/SB2/n2645 ), .C(\U1/aes_core/SB2/n2644 ), .D(
        \U1/aes_core/SB2/n2945 ), .Y(\U1/aes_core/SB2/n2653 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U302  ( .A0(\U1/aes_core/SB2/n2647 ), 
        .A1(\U1/aes_core/SB2/n2912 ), .B0(\U1/aes_core/SB2/n2809 ), .Y(
        \U1/aes_core/SB2/n2649 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U299  ( .A(\U1/aes_core/SB2/n2865 ), .B(
        \U1/aes_core/SB2/n2933 ), .Y(\U1/aes_core/SB2/n2876 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U298  ( .A0(\U1/aes_core/SB2/n2755 ), 
        .A1(\U1/aes_core/SB2/n2955 ), .B0(\U1/aes_core/SB2/n2876 ), .B1(
        \U1/aes_core/SB2/n2908 ), .C0(\U1/aes_core/SB2/n2949 ), .C1(
        \U1/aes_core/SB2/n2958 ), .Y(\U1/aes_core/SB2/n2651 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U297  ( .A(\U1/aes_core/SB2/n2656 ), .B(
        \U1/aes_core/SB2/n2655 ), .C(\U1/aes_core/SB2/n2654 ), .D(
        \U1/aes_core/SB2/n2653 ), .E(\U1/aes_core/SB2/n2652 ), .F(
        \U1/aes_core/SB2/n2651 ), .Y(\U1/aes_core/SB2/n2839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U296  ( .AN(\U1/aes_core/SB2/n2660 ), 
        .B(\U1/aes_core/SB2/n2659 ), .C(\U1/aes_core/SB2/n2658 ), .D(
        \U1/aes_core/SB2/n2657 ), .Y(\U1/aes_core/SB2/n2670 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U295  ( .A0(\U1/aes_core/SB2/n2943 ), 
        .A1(\U1/aes_core/SB2/n2832 ), .B0(\U1/aes_core/SB2/n2938 ), .B1(
        \U1/aes_core/SB2/n2831 ), .C0(\U1/aes_core/SB2/n2661 ), .C1(
        \U1/aes_core/SB2/n2953 ), .Y(\U1/aes_core/SB2/n2669 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U294  ( .A0(\U1/aes_core/SB2/n2907 ), 
        .A1(\U1/aes_core/SB2/n2792 ), .B0(\U1/aes_core/SB2/n2662 ), .B1(
        \U1/aes_core/SB2/n2755 ), .Y(\U1/aes_core/SB2/n2663 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U293  ( .A0(\U1/aes_core/SB2/n2809 ), 
        .A1(\U1/aes_core/SB2/n2826 ), .B0(\U1/aes_core/SB2/n2825 ), .B1(
        \U1/aes_core/SB2/n2910 ), .C0(\U1/aes_core/SB2/n2663 ), .Y(
        \U1/aes_core/SB2/n2668 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U292  ( .A(\U1/aes_core/SB2/n2918 ), .B(
        \U1/aes_core/SB2/n2957 ), .Y(\U1/aes_core/SB2/n2665 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U291  ( .A0(\U1/aes_core/SB2/n2747 ), 
        .A1(\U1/aes_core/SB2/n2666 ), .B0(\U1/aes_core/SB2/n2939 ), .B1(
        \U1/aes_core/SB2/n2665 ), .C0(\U1/aes_core/SB2/n2664 ), .Y(
        \U1/aes_core/SB2/n2667 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U290  ( .AN(\U1/aes_core/SB2/n2670 ), 
        .B(\U1/aes_core/SB2/n2669 ), .C(\U1/aes_core/SB2/n2668 ), .D(
        \U1/aes_core/SB2/n2667 ), .Y(\U1/aes_core/SB2/n2884 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U289  ( .A(\U1/aes_core/SB2/n2671 ), .Y(
        \U1/aes_core/SB2/n2687 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U288  ( .A0(\U1/aes_core/SB2/n2776 ), 
        .A1(\U1/aes_core/SB2/n2845 ), .B0(\U1/aes_core/SB2/n2672 ), .Y(
        \U1/aes_core/SB2/n2686 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U287  ( .A0(\U1/aes_core/SB2/n2939 ), 
        .A1(\U1/aes_core/SB2/n2938 ), .B0(\U1/aes_core/SB2/n2909 ), .B1(
        \U1/aes_core/SB2/n2673 ), .Y(\U1/aes_core/SB2/n2674 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U286  ( .A0(\U1/aes_core/SB2/n2920 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2936 ), .B1(
        \U1/aes_core/SB2/n2948 ), .C0(\U1/aes_core/SB2/n2674 ), .Y(
        \U1/aes_core/SB2/n2685 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U285  ( .A(\U1/aes_core/SB2/n2678 ), .B(
        \U1/aes_core/SB2/n2677 ), .C(\U1/aes_core/SB2/n2676 ), .D(
        \U1/aes_core/SB2/n2675 ), .Y(\U1/aes_core/SB2/n2684 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U284  ( .AN(\U1/aes_core/SB2/n2682 ), 
        .B(\U1/aes_core/SB2/n2681 ), .C(\U1/aes_core/SB2/n2680 ), .D(
        \U1/aes_core/SB2/n2679 ), .Y(\U1/aes_core/SB2/n2683 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U283  ( .A(\U1/aes_core/SB2/n2688 ), .B(
        \U1/aes_core/SB2/n2687 ), .C(\U1/aes_core/SB2/n2686 ), .D(
        \U1/aes_core/SB2/n2685 ), .E(\U1/aes_core/SB2/n2684 ), .F(
        \U1/aes_core/SB2/n2683 ), .Y(\U1/aes_core/SB2/n2788 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U282  ( .A0(\U1/aes_core/SB2/n2875 ), 
        .A1(\U1/aes_core/SB2/n2792 ), .B0(\U1/aes_core/SB2/n2689 ), .Y(
        \U1/aes_core/SB2/n2704 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U281  ( .AN(\U1/aes_core/SB2/n2693 ), 
        .B(\U1/aes_core/SB2/n2692 ), .C(\U1/aes_core/SB2/n2691 ), .D(
        \U1/aes_core/SB2/n2690 ), .Y(\U1/aes_core/SB2/n2703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U280  ( .A(\U1/aes_core/SB2/n2930 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2944 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U279  ( .A(\U1/aes_core/SB2/n2696 ), .B(
        \U1/aes_core/SB2/n2695 ), .C(\U1/aes_core/SB2/n2694 ), .D(
        \U1/aes_core/SB2/n2944 ), .Y(\U1/aes_core/SB2/n2702 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U278  ( .A(\U1/aes_core/SB2/n2700 ), .B(
        \U1/aes_core/SB2/n2699 ), .C(\U1/aes_core/SB2/n2698 ), .D(
        \U1/aes_core/SB2/n2697 ), .Y(\U1/aes_core/SB2/n2701 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U277  ( .A(\U1/aes_core/SB2/n2706 ), .B(
        \U1/aes_core/SB2/n2705 ), .C(\U1/aes_core/SB2/n2704 ), .D(
        \U1/aes_core/SB2/n2703 ), .E(\U1/aes_core/SB2/n2702 ), .F(
        \U1/aes_core/SB2/n2701 ), .Y(\U1/aes_core/SB2/n2812 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U276  ( .AN(\U1/aes_core/SB2/n2710 ), 
        .B(\U1/aes_core/SB2/n2709 ), .C(\U1/aes_core/SB2/n2708 ), .D(
        \U1/aes_core/SB2/n2707 ), .Y(\U1/aes_core/SB2/n2719 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U275  ( .A(\U1/aes_core/SB2/n2714 ), .B(
        \U1/aes_core/SB2/n2713 ), .C(\U1/aes_core/SB2/n2712 ), .D(
        \U1/aes_core/SB2/n2711 ), .Y(\U1/aes_core/SB2/n2718 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U274  ( .A(\U1/aes_core/SB2/n2874 ), .B(
        \U1/aes_core/SB2/n2931 ), .C(\U1/aes_core/SB2/n2933 ), .Y(
        \U1/aes_core/SB2/n2716 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U273  ( .A0(\U1/aes_core/SB2/n2716 ), 
        .A1(\U1/aes_core/SB2/n2921 ), .B0(\U1/aes_core/SB2/n2755 ), .B1(
        \U1/aes_core/SB2/n2957 ), .C0(\U1/aes_core/SB2/n2715 ), .Y(
        \U1/aes_core/SB2/n2717 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U272  ( .A(\U1/aes_core/SB2/n2722 ), .B(
        \U1/aes_core/SB2/n2721 ), .C(\U1/aes_core/SB2/n2720 ), .D(
        \U1/aes_core/SB2/n2719 ), .E(\U1/aes_core/SB2/n2718 ), .F(
        \U1/aes_core/SB2/n2717 ), .Y(\U1/aes_core/SB2/n2860 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U271  ( .A0(\U1/aes_core/SB2/n2755 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2723 ), .Y(
        \U1/aes_core/SB2/n2737 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U270  ( .A0(\U1/aes_core/SB2/n2864 ), 
        .A1(\U1/aes_core/SB2/n2866 ), .B0(\U1/aes_core/SB2/n2942 ), .B1(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2724 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U269  ( .A0(\U1/aes_core/SB2/n2775 ), 
        .A1(\U1/aes_core/SB2/n2863 ), .B0(\U1/aes_core/SB2/n2776 ), .B1(
        \U1/aes_core/SB2/n2840 ), .C0(\U1/aes_core/SB2/n2724 ), .Y(
        \U1/aes_core/SB2/n2736 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U268  ( .A(\U1/aes_core/SB2/n2725 ), .Y(
        \U1/aes_core/SB2/n2728 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U267  ( .AN(\U1/aes_core/SB2/n2729 ), 
        .B(\U1/aes_core/SB2/n2728 ), .C(\U1/aes_core/SB2/n2727 ), .D(
        \U1/aes_core/SB2/n2726 ), .Y(\U1/aes_core/SB2/n2735 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U266  ( .A(\U1/aes_core/SB2/n2733 ), .B(
        \U1/aes_core/SB2/n2732 ), .C(\U1/aes_core/SB2/n2731 ), .D(
        \U1/aes_core/SB2/n2730 ), .Y(\U1/aes_core/SB2/n2734 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U265  ( .A(\U1/aes_core/SB2/n2739 ), .B(
        \U1/aes_core/SB2/n2738 ), .C(\U1/aes_core/SB2/n2737 ), .D(
        \U1/aes_core/SB2/n2736 ), .E(\U1/aes_core/SB2/n2735 ), .F(
        \U1/aes_core/SB2/n2734 ), .Y(\U1/aes_core/SB2/n2819 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U264  ( .A0(\U1/aes_core/SB2/n2931 ), 
        .A1(\U1/aes_core/SB2/n2740 ), .B0(\U1/aes_core/SB2/n2941 ), .B1(
        \U1/aes_core/SB2/n2866 ), .Y(\U1/aes_core/SB2/n2741 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U263  ( .A0(\U1/aes_core/SB2/n2792 ), 
        .A1(\U1/aes_core/SB2/n2958 ), .B0(\U1/aes_core/SB2/n2742 ), .B1(
        \U1/aes_core/SB2/n2948 ), .C0(\U1/aes_core/SB2/n2741 ), .Y(
        \U1/aes_core/SB2/n2754 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U262  ( .AN(\U1/aes_core/SB2/n2746 ), 
        .B(\U1/aes_core/SB2/n2745 ), .C(\U1/aes_core/SB2/n2744 ), .D(
        \U1/aes_core/SB2/n2743 ), .Y(\U1/aes_core/SB2/n2753 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U261  ( .A0(\U1/aes_core/SB2/n2951 ), 
        .A1(\U1/aes_core/SB2/n2747 ), .B0(\U1/aes_core/SB2/n2942 ), .Y(
        \U1/aes_core/SB2/n2751 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U260  ( .A(\U1/aes_core/SB2/n2918 ), .B(
        \U1/aes_core/SB2/n2923 ), .Y(\U1/aes_core/SB2/n2748 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U259  ( .A0(\U1/aes_core/SB2/n2873 ), 
        .A1(\U1/aes_core/SB2/n2748 ), .B0(\U1/aes_core/SB2/n2874 ), .B1(
        \U1/aes_core/SB2/n2820 ), .Y(\U1/aes_core/SB2/n2749 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U258  ( .A(\U1/aes_core/SB2/n2751 ), .B(
        \U1/aes_core/SB2/n2750 ), .C(\U1/aes_core/SB2/n2749 ), .Y(
        \U1/aes_core/SB2/n2752 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U257  ( .A(\U1/aes_core/SB2/n2812 ), .B(
        \U1/aes_core/SB2/n2860 ), .C(\U1/aes_core/SB2/n2819 ), .D(
        \U1/aes_core/SB2/n2754 ), .E(\U1/aes_core/SB2/n2753 ), .F(
        \U1/aes_core/SB2/n2752 ), .Y(\U1/aes_core/SB2/n2927 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U256  ( .A(\U1/aes_core/SB2/n2839 ), .B(
        \U1/aes_core/SB2/n2884 ), .C(\U1/aes_core/SB2/n2788 ), .D(
        \U1/aes_core/SB2/n2927 ), .Y(\U1/aes_core/SB2/n2768 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U255  ( .A0(\U1/aes_core/SB2/n2907 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2755 ), .B1(
        \U1/aes_core/SB2/n2923 ), .Y(\U1/aes_core/SB2/n2756 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U254  ( .A0(\U1/aes_core/SB2/n2912 ), 
        .A1(\U1/aes_core/SB2/n2930 ), .B0(\U1/aes_core/SB2/n2943 ), .B1(
        \U1/aes_core/SB2/n2951 ), .C0(\U1/aes_core/SB2/n2756 ), .Y(
        \U1/aes_core/SB2/n2767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U253  ( .A(\U1/aes_core/SB2/n2757 ), .Y(
        \U1/aes_core/SB2/n2760 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U252  ( .A0(\U1/aes_core/SB2/n2758 ), 
        .A1(\U1/aes_core/SB2/n2863 ), .B0(\U1/aes_core/SB2/n2791 ), .B1(
        \U1/aes_core/SB2/n2843 ), .Y(\U1/aes_core/SB2/n2759 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U251  ( .A0(\U1/aes_core/SB2/n2931 ), 
        .A1(\U1/aes_core/SB2/n2760 ), .B0(\U1/aes_core/SB2/n2913 ), .B1(
        \U1/aes_core/SB2/n2841 ), .C0(\U1/aes_core/SB2/n2759 ), .Y(
        \U1/aes_core/SB2/n2766 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U250  ( .A0(\U1/aes_core/SB2/n2953 ), 
        .A1(\U1/aes_core/SB2/n2809 ), .B0(\U1/aes_core/SB2/n2933 ), .Y(
        \U1/aes_core/SB2/n2764 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB2/U249  ( .A(\U1/aes_core/SB2/n2764 ), .B(
        \U1/aes_core/SB2/n2763 ), .C(\U1/aes_core/SB2/n2762 ), .D(
        \U1/aes_core/SB2/n2761 ), .Y(\U1/aes_core/SB2/n2765 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U248  ( .AN(\U1/aes_core/SB2/n2768 ), 
        .B(\U1/aes_core/SB2/n2767 ), .C(\U1/aes_core/SB2/n2766 ), .D(
        \U1/aes_core/SB2/n2765 ), .Y(\U1/aes_core/sb2 [27]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U247  ( .A0(\U1/aes_core/SB2/n2783 ), 
        .A1(\U1/aes_core/SB2/n2919 ), .B0(\U1/aes_core/SB2/n2842 ), .Y(
        \U1/aes_core/SB2/n2780 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U246  ( .A(\U1/aes_core/SB2/n2771 ), .B(
        \U1/aes_core/SB2/n2770 ), .C(\U1/aes_core/SB2/n2769 ), .Y(
        \U1/aes_core/SB2/n2779 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U245  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2942 ), .Y(\U1/aes_core/SB2/n2774 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U244  ( .A(\U1/aes_core/SB2/n2913 ), .B(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2772 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U243  ( .A0(\U1/aes_core/SB2/n2774 ), 
        .A1(\U1/aes_core/SB2/n2773 ), .B0(\U1/aes_core/SB2/n2772 ), .B1(
        \U1/aes_core/SB2/n2936 ), .C0(\U1/aes_core/SB2/n2919 ), .C1(
        \U1/aes_core/SB2/n2824 ), .Y(\U1/aes_core/SB2/n2778 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U242  ( .A0(\U1/aes_core/SB2/n2875 ), 
        .A1(\U1/aes_core/SB2/n2776 ), .B0(\U1/aes_core/SB2/n2958 ), .B1(
        \U1/aes_core/SB2/n2948 ), .C0(\U1/aes_core/SB2/n2921 ), .C1(
        \U1/aes_core/SB2/n2775 ), .Y(\U1/aes_core/SB2/n2777 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U241  ( .A(\U1/aes_core/SB2/n2782 ), .B(
        \U1/aes_core/SB2/n2781 ), .C(\U1/aes_core/SB2/n2780 ), .D(
        \U1/aes_core/SB2/n2779 ), .E(\U1/aes_core/SB2/n2778 ), .F(
        \U1/aes_core/SB2/n2777 ), .Y(\U1/aes_core/SB2/n2928 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U240  ( .A0(\U1/aes_core/SB2/n2783 ), 
        .A1(\U1/aes_core/SB2/n2792 ), .B0(\U1/aes_core/SB2/n2863 ), .Y(
        \U1/aes_core/SB2/n2818 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB2/U239  ( .A0(\U1/aes_core/SB2/n2908 ), 
        .A1(\U1/aes_core/SB2/n2921 ), .A2(\U1/aes_core/SB2/n2840 ), .B0(
        \U1/aes_core/SB2/n2937 ), .Y(\U1/aes_core/SB2/n2817 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U238  ( .A(\U1/aes_core/SB2/n2787 ), .B(
        \U1/aes_core/SB2/n2786 ), .C(\U1/aes_core/SB2/n2785 ), .D(
        \U1/aes_core/SB2/n2784 ), .Y(\U1/aes_core/SB2/n2814 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U237  ( .A(\U1/aes_core/SB2/n2788 ), .Y(
        \U1/aes_core/SB2/n2811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U236  ( .A(\U1/aes_core/SB2/n2789 ), .Y(
        \U1/aes_core/SB2/n2805 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB2/U235  ( .A0(\U1/aes_core/SB2/n2791 ), 
        .A1(\U1/aes_core/SB2/n2949 ), .B0N(\U1/aes_core/SB2/n2790 ), .Y(
        \U1/aes_core/SB2/n2804 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U234  ( .A0(\U1/aes_core/SB2/n2956 ), 
        .A1(\U1/aes_core/SB2/n2792 ), .B0(\U1/aes_core/SB2/n2842 ), .B1(
        \U1/aes_core/SB2/n2923 ), .C0(\U1/aes_core/SB2/n2937 ), .C1(
        \U1/aes_core/SB2/n2958 ), .Y(\U1/aes_core/SB2/n2803 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U233  ( .AN(\U1/aes_core/SB2/n2796 ), 
        .B(\U1/aes_core/SB2/n2795 ), .C(\U1/aes_core/SB2/n2794 ), .D(
        \U1/aes_core/SB2/n2793 ), .Y(\U1/aes_core/SB2/n2802 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U232  ( .A(\U1/aes_core/SB2/n2800 ), .B(
        \U1/aes_core/SB2/n2799 ), .C(\U1/aes_core/SB2/n2798 ), .D(
        \U1/aes_core/SB2/n2797 ), .Y(\U1/aes_core/SB2/n2801 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U231  ( .A(\U1/aes_core/SB2/n2806 ), .B(
        \U1/aes_core/SB2/n2805 ), .C(\U1/aes_core/SB2/n2804 ), .D(
        \U1/aes_core/SB2/n2803 ), .E(\U1/aes_core/SB2/n2802 ), .F(
        \U1/aes_core/SB2/n2801 ), .Y(\U1/aes_core/SB2/n2807 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U230  ( .A(\U1/aes_core/SB2/n2807 ), .Y(
        \U1/aes_core/SB2/n2906 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U229  ( .A0(\U1/aes_core/SB2/n2875 ), 
        .A1(\U1/aes_core/SB2/n2918 ), .B0(\U1/aes_core/SB2/n2958 ), .B1(
        \U1/aes_core/SB2/n2957 ), .Y(\U1/aes_core/SB2/n2808 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U228  ( .A0(\U1/aes_core/SB2/n2865 ), 
        .A1(\U1/aes_core/SB2/n2809 ), .B0(\U1/aes_core/SB2/n2910 ), .B1(
        \U1/aes_core/SB2/n2932 ), .C0(\U1/aes_core/SB2/n2808 ), .Y(
        \U1/aes_core/SB2/n2810 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U227  ( .AN(\U1/aes_core/SB2/n2812 ), 
        .B(\U1/aes_core/SB2/n2811 ), .C(\U1/aes_core/SB2/n2906 ), .D(
        \U1/aes_core/SB2/n2810 ), .Y(\U1/aes_core/SB2/n2813 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U226  ( .A(\U1/aes_core/SB2/n2818 ), .B(
        \U1/aes_core/SB2/n2817 ), .C(\U1/aes_core/SB2/n2816 ), .D(
        \U1/aes_core/SB2/n2815 ), .E(\U1/aes_core/SB2/n2814 ), .F(
        \U1/aes_core/SB2/n2813 ), .Y(\U1/aes_core/SB2/n2883 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U225  ( .A(\U1/aes_core/SB2/n2819 ), .Y(
        \U1/aes_core/SB2/n2823 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U224  ( .A0(\U1/aes_core/SB2/n2821 ), 
        .A1(\U1/aes_core/SB2/n2820 ), .B0(\U1/aes_core/SB2/n2867 ), .B1(
        \U1/aes_core/SB2/n2826 ), .Y(\U1/aes_core/SB2/n2822 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U223  ( .A0(\U1/aes_core/SB2/n2937 ), 
        .A1(\U1/aes_core/SB2/n2824 ), .B0(\U1/aes_core/SB2/n2823 ), .C0(
        \U1/aes_core/SB2/n2822 ), .Y(\U1/aes_core/SB2/n2838 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U222  ( .A0(\U1/aes_core/SB2/n2825 ), 
        .A1(\U1/aes_core/SB2/n2909 ), .B0(\U1/aes_core/SB2/n2938 ), .Y(
        \U1/aes_core/SB2/n2830 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U221  ( .A0(\U1/aes_core/SB2/n2826 ), 
        .A1(\U1/aes_core/SB2/n2912 ), .B0(\U1/aes_core/SB2/n2941 ), .Y(
        \U1/aes_core/SB2/n2829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U220  ( .A(\U1/aes_core/SB2/n2830 ), .B(
        \U1/aes_core/SB2/n2829 ), .C(\U1/aes_core/SB2/n2828 ), .D(
        \U1/aes_core/SB2/n2827 ), .Y(\U1/aes_core/SB2/n2837 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U219  ( .A(\U1/aes_core/SB2/n2868 ), .B(
        \U1/aes_core/SB2/n2831 ), .Y(\U1/aes_core/SB2/n2835 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U218  ( .A(\U1/aes_core/SB2/n2832 ), .B(
        \U1/aes_core/SB2/n2873 ), .Y(\U1/aes_core/SB2/n2834 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U217  ( .A0(\U1/aes_core/SB2/n2835 ), 
        .A1(\U1/aes_core/SB2/n2955 ), .B0(\U1/aes_core/SB2/n2834 ), .B1(
        \U1/aes_core/SB2/n2919 ), .C0(\U1/aes_core/SB2/n2833 ), .C1(
        \U1/aes_core/SB2/n2920 ), .Y(\U1/aes_core/SB2/n2836 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U216  ( .A(\U1/aes_core/SB2/n2928 ), .B(
        \U1/aes_core/SB2/n2883 ), .C(\U1/aes_core/SB2/n2839 ), .D(
        \U1/aes_core/SB2/n2838 ), .E(\U1/aes_core/SB2/n2837 ), .F(
        \U1/aes_core/SB2/n2836 ), .Y(\U1/aes_core/sb2 [28]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U215  ( .A1N(\U1/aes_core/SB2/n2841 ), 
        .A0(\U1/aes_core/SB2/n2840 ), .B0(\U1/aes_core/SB2/n2918 ), .Y(
        \U1/aes_core/SB2/n2857 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U214  ( .A(\U1/aes_core/SB2/n2931 ), .B(
        \U1/aes_core/SB2/n2912 ), .Y(\U1/aes_core/SB2/n2844 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U213  ( .A0(\U1/aes_core/SB2/n2955 ), 
        .A1(\U1/aes_core/SB2/n2845 ), .B0(\U1/aes_core/SB2/n2844 ), .B1(
        \U1/aes_core/SB2/n2958 ), .C0(\U1/aes_core/SB2/n2843 ), .C1(
        \U1/aes_core/SB2/n2842 ), .Y(\U1/aes_core/SB2/n2856 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U212  ( .A(\U1/aes_core/SB2/n2846 ), .Y(
        \U1/aes_core/SB2/n2849 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U211  ( .AN(\U1/aes_core/SB2/n2850 ), 
        .B(\U1/aes_core/SB2/n2849 ), .C(\U1/aes_core/SB2/n2848 ), .D(
        \U1/aes_core/SB2/n2847 ), .Y(\U1/aes_core/SB2/n2855 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U210  ( .A(\U1/aes_core/SB2/n2853 ), .B(
        \U1/aes_core/SB2/n2852 ), .C(\U1/aes_core/SB2/n2851 ), .Y(
        \U1/aes_core/SB2/n2854 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U209  ( .A(\U1/aes_core/SB2/n2859 ), .B(
        \U1/aes_core/SB2/n2858 ), .C(\U1/aes_core/SB2/n2857 ), .D(
        \U1/aes_core/SB2/n2856 ), .E(\U1/aes_core/SB2/n2855 ), .F(
        \U1/aes_core/SB2/n2854 ), .Y(\U1/aes_core/SB2/n2929 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U208  ( .A(\U1/aes_core/SB2/n2860 ), .Y(
        \U1/aes_core/SB2/n2862 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U207  ( .A0(\U1/aes_core/SB2/n2942 ), 
        .A1(\U1/aes_core/SB2/n2939 ), .B0(\U1/aes_core/SB2/n2943 ), .B1(
        \U1/aes_core/SB2/n2941 ), .Y(\U1/aes_core/SB2/n2861 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U206  ( .A0(\U1/aes_core/SB2/n2918 ), 
        .A1(\U1/aes_core/SB2/n2863 ), .B0(\U1/aes_core/SB2/n2862 ), .C0(
        \U1/aes_core/SB2/n2861 ), .Y(\U1/aes_core/SB2/n2882 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U205  ( .A0(\U1/aes_core/SB2/n2865 ), 
        .A1(\U1/aes_core/SB2/n2942 ), .B0(\U1/aes_core/SB2/n2864 ), .Y(
        \U1/aes_core/SB2/n2871 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U204  ( .A0(\U1/aes_core/SB2/n2868 ), 
        .A1(\U1/aes_core/SB2/n2867 ), .B0(\U1/aes_core/SB2/n2866 ), .Y(
        \U1/aes_core/SB2/n2870 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U203  ( .AN(\U1/aes_core/SB2/n2872 ), 
        .B(\U1/aes_core/SB2/n2871 ), .C(\U1/aes_core/SB2/n2870 ), .D(
        \U1/aes_core/SB2/n2869 ), .Y(\U1/aes_core/SB2/n2881 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U202  ( .A0(\U1/aes_core/SB2/n2938 ), 
        .A1(\U1/aes_core/SB2/n2874 ), .B0(\U1/aes_core/SB2/n2873 ), .Y(
        \U1/aes_core/SB2/n2878 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB2/U201  ( .A0(\U1/aes_core/SB2/n2920 ), .A1(
        \U1/aes_core/SB2/n2876 ), .B0(\U1/aes_core/SB2/n2957 ), .B1(
        \U1/aes_core/SB2/n2875 ), .Y(\U1/aes_core/SB2/n2877 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U200  ( .A0(\U1/aes_core/SB2/n2879 ), 
        .A1(\U1/aes_core/SB2/n2919 ), .B0(\U1/aes_core/SB2/n2878 ), .C0(
        \U1/aes_core/SB2/n2877 ), .Y(\U1/aes_core/SB2/n2880 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U199  ( .A(\U1/aes_core/SB2/n2929 ), .B(
        \U1/aes_core/SB2/n2884 ), .C(\U1/aes_core/SB2/n2883 ), .D(
        \U1/aes_core/SB2/n2882 ), .E(\U1/aes_core/SB2/n2881 ), .F(
        \U1/aes_core/SB2/n2880 ), .Y(\U1/aes_core/sb2 [29]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U198  ( .A0(\U1/aes_core/SB2/n3212 ), 
        .A1(\U1/aes_core/SB2/n3232 ), .B0(\U1/aes_core/SB2/n3253 ), .B1(
        \U1/aes_core/SB2/n3243 ), .Y(\U1/aes_core/SB2/n2885 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U197  ( .A0(\U1/aes_core/SB2/n3163 ), 
        .A1(\U1/aes_core/SB2/n3257 ), .B0(\U1/aes_core/SB2/n3113 ), .B1(
        \U1/aes_core/SB2/n3184 ), .C0(\U1/aes_core/SB2/n2885 ), .Y(
        \U1/aes_core/SB2/n2891 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U196  ( .A(\U1/aes_core/SB2/n3238 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3047 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U195  ( .A(\U1/aes_core/SB2/n3212 ), .B(
        \U1/aes_core/SB2/n3188 ), .Y(\U1/aes_core/SB2/n3028 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U194  ( .A(\U1/aes_core/SB2/n3232 ), .B(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n2996 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U193  ( .A(\U1/aes_core/SB2/n3152 ), .B(
        \U1/aes_core/SB2/n3195 ), .Y(\U1/aes_core/SB2/n3015 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U192  ( .A(\U1/aes_core/SB2/n3047 ), .B(
        \U1/aes_core/SB2/n3028 ), .C(\U1/aes_core/SB2/n2996 ), .D(
        \U1/aes_core/SB2/n3015 ), .Y(\U1/aes_core/SB2/n2890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U191  ( .A(\U1/aes_core/SB2/n3258 ), .B(
        \U1/aes_core/SB2/n3236 ), .Y(\U1/aes_core/SB2/n3141 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U190  ( .A0(\U1/aes_core/SB2/n3189 ), 
        .A1(\U1/aes_core/SB2/n3141 ), .B0(\U1/aes_core/SB2/n3242 ), .Y(
        \U1/aes_core/SB2/n2888 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U189  ( .A0(\U1/aes_core/SB2/n3239 ), 
        .A1(\U1/aes_core/SB2/n3130 ), .B0(\U1/aes_core/SB2/n3142 ), .Y(
        \U1/aes_core/SB2/n2887 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U188  ( .A0(\U1/aes_core/SB2/n3147 ), 
        .A1(\U1/aes_core/SB2/n3187 ), .B0(\U1/aes_core/SB2/n3241 ), .Y(
        \U1/aes_core/SB2/n2886 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U187  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3239 ), .Y(\U1/aes_core/SB2/n3114 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U186  ( .A(\U1/aes_core/SB2/n2888 ), .B(
        \U1/aes_core/SB2/n2887 ), .C(\U1/aes_core/SB2/n2886 ), .D(
        \U1/aes_core/SB2/n3114 ), .Y(\U1/aes_core/SB2/n2889 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U185  ( .A(\U1/aes_core/SB2/n2894 ), .B(
        \U1/aes_core/SB2/n2893 ), .C(\U1/aes_core/SB2/n2892 ), .D(
        \U1/aes_core/SB2/n2891 ), .E(\U1/aes_core/SB2/n2890 ), .F(
        \U1/aes_core/SB2/n2889 ), .Y(\U1/aes_core/SB2/n3262 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U184  ( .A0(\U1/aes_core/SB2/n3068 ), 
        .A1(\U1/aes_core/SB2/n3243 ), .B0(\U1/aes_core/SB2/n3251 ), .B1(
        \U1/aes_core/SB2/n3186 ), .C0(\U1/aes_core/SB2/n3262 ), .Y(
        \U1/aes_core/SB2/n2895 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U183  ( .A(\U1/aes_core/SB2/n2895 ), .Y(
        \U1/aes_core/SB2/n2902 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U182  ( .A(\U1/aes_core/SB2/n3195 ), .B(
        \U1/aes_core/SB2/n2982 ), .Y(\U1/aes_core/SB2/n3104 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U181  ( .A1N(\U1/aes_core/SB2/n3104 ), 
        .A0(\U1/aes_core/SB2/n3213 ), .B0(\U1/aes_core/SB2/n3185 ), .Y(
        \U1/aes_core/SB2/n2898 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U180  ( .A0(\U1/aes_core/SB2/n3153 ), 
        .A1(\U1/aes_core/SB2/n3061 ), .B0(\U1/aes_core/SB2/n3212 ), .Y(
        \U1/aes_core/SB2/n2897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U179  ( .A0(\U1/aes_core/SB2/n3239 ), 
        .A1(\U1/aes_core/SB2/n3194 ), .B0(\U1/aes_core/SB2/n3233 ), .Y(
        \U1/aes_core/SB2/n2896 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U178  ( .A(\U1/aes_core/SB2/n3210 ), .B(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n3011 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U177  ( .A(\U1/aes_core/SB2/n2898 ), .B(
        \U1/aes_core/SB2/n2897 ), .C(\U1/aes_core/SB2/n2896 ), .D(
        \U1/aes_core/SB2/n3011 ), .Y(\U1/aes_core/SB2/n2901 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U176  ( .A(\U1/aes_core/SB2/n3209 ), .B(
        \U1/aes_core/SB2/n3241 ), .Y(\U1/aes_core/SB2/n3240 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U175  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3187 ), .Y(\U1/aes_core/SB2/n2899 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U174  ( .A0(\U1/aes_core/SB2/n3240 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n2899 ), .B1(
        \U1/aes_core/SB2/n3221 ), .C0(\U1/aes_core/SB2/n3164 ), .C1(
        \U1/aes_core/SB2/n3166 ), .Y(\U1/aes_core/SB2/n2900 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U173  ( .A(\U1/aes_core/SB2/n2905 ), .B(
        \U1/aes_core/SB2/n2904 ), .C(\U1/aes_core/SB2/n2903 ), .D(
        \U1/aes_core/SB2/n2902 ), .E(\U1/aes_core/SB2/n2901 ), .F(
        \U1/aes_core/SB2/n2900 ), .Y(\U1/aes_core/sb2 [2]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U172  ( .A0(\U1/aes_core/SB2/n2908 ), 
        .A1(\U1/aes_core/SB2/n2948 ), .B0(\U1/aes_core/SB2/n2907 ), .B1(
        \U1/aes_core/SB2/n2955 ), .C0(\U1/aes_core/SB2/n2906 ), .Y(
        \U1/aes_core/SB2/n2926 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U171  ( .A0(\U1/aes_core/SB2/n2909 ), 
        .A1(\U1/aes_core/SB2/n2953 ), .B0(\U1/aes_core/SB2/n2942 ), .Y(
        \U1/aes_core/SB2/n2917 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U170  ( .A0(\U1/aes_core/SB2/n2933 ), 
        .A1(\U1/aes_core/SB2/n2910 ), .B0(\U1/aes_core/SB2/n2941 ), .Y(
        \U1/aes_core/SB2/n2916 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U169  ( .A0(\U1/aes_core/SB2/n2913 ), 
        .A1(\U1/aes_core/SB2/n2912 ), .B0(\U1/aes_core/SB2/n2911 ), .Y(
        \U1/aes_core/SB2/n2915 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U168  ( .A(\U1/aes_core/SB2/n2917 ), .B(
        \U1/aes_core/SB2/n2916 ), .C(\U1/aes_core/SB2/n2915 ), .D(
        \U1/aes_core/SB2/n2914 ), .Y(\U1/aes_core/SB2/n2925 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U167  ( .A(\U1/aes_core/SB2/n2948 ), .B(
        \U1/aes_core/SB2/n2918 ), .Y(\U1/aes_core/SB2/n2950 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U166  ( .A(\U1/aes_core/SB2/n2938 ), .B(
        \U1/aes_core/SB2/n2950 ), .Y(\U1/aes_core/SB2/n2922 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U165  ( .A0(\U1/aes_core/SB2/n2936 ), 
        .A1(\U1/aes_core/SB2/n2923 ), .B0(\U1/aes_core/SB2/n2922 ), .B1(
        \U1/aes_core/SB2/n2921 ), .C0(\U1/aes_core/SB2/n2920 ), .C1(
        \U1/aes_core/SB2/n2919 ), .Y(\U1/aes_core/SB2/n2924 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U164  ( .A(\U1/aes_core/SB2/n2929 ), .B(
        \U1/aes_core/SB2/n2928 ), .C(\U1/aes_core/SB2/n2927 ), .D(
        \U1/aes_core/SB2/n2926 ), .E(\U1/aes_core/SB2/n2925 ), .F(
        \U1/aes_core/SB2/n2924 ), .Y(\U1/aes_core/sb2 [30]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U163  ( .A0(\U1/aes_core/SB2/n2933 ), 
        .A1(\U1/aes_core/SB2/n2932 ), .B0(\U1/aes_core/SB2/n2931 ), .B1(
        \U1/aes_core/SB2/n2930 ), .Y(\U1/aes_core/SB2/n2934 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U162  ( .A0(\U1/aes_core/SB2/n2937 ), 
        .A1(\U1/aes_core/SB2/n2936 ), .B0(\U1/aes_core/SB2/n2935 ), .C0(
        \U1/aes_core/SB2/n2934 ), .Y(\U1/aes_core/SB2/n2961 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U161  ( .A1N(\U1/aes_core/SB2/n2940 ), 
        .A0(\U1/aes_core/SB2/n2939 ), .B0(\U1/aes_core/SB2/n2938 ), .Y(
        \U1/aes_core/SB2/n2947 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U160  ( .A0(\U1/aes_core/SB2/n2943 ), 
        .A1(\U1/aes_core/SB2/n2942 ), .B0(\U1/aes_core/SB2/n2941 ), .Y(
        \U1/aes_core/SB2/n2946 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U159  ( .A(\U1/aes_core/SB2/n2947 ), .B(
        \U1/aes_core/SB2/n2946 ), .C(\U1/aes_core/SB2/n2945 ), .D(
        \U1/aes_core/SB2/n2944 ), .Y(\U1/aes_core/SB2/n2960 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U158  ( .A(\U1/aes_core/SB2/n2949 ), .B(
        \U1/aes_core/SB2/n2948 ), .Y(\U1/aes_core/SB2/n2952 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U157  ( .A0(\U1/aes_core/SB2/n2953 ), 
        .A1(\U1/aes_core/SB2/n2952 ), .B0(\U1/aes_core/SB2/n2951 ), .B1(
        \U1/aes_core/SB2/n2950 ), .Y(\U1/aes_core/SB2/n2954 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U156  ( .A0(\U1/aes_core/SB2/n2958 ), 
        .A1(\U1/aes_core/SB2/n2957 ), .B0(\U1/aes_core/SB2/n2956 ), .B1(
        \U1/aes_core/SB2/n2955 ), .C0(\U1/aes_core/SB2/n2954 ), .Y(
        \U1/aes_core/SB2/n2959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U155  ( .A(\U1/aes_core/SB2/n2964 ), .B(
        \U1/aes_core/SB2/n2963 ), .C(\U1/aes_core/SB2/n2962 ), .D(
        \U1/aes_core/SB2/n2961 ), .E(\U1/aes_core/SB2/n2960 ), .F(
        \U1/aes_core/SB2/n2959 ), .Y(\U1/aes_core/sb2 [31]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U154  ( .A(\U1/aes_core/SB2/n3068 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3245 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U153  ( .AN(\U1/aes_core/SB2/n2967 ), 
        .B(\U1/aes_core/SB2/n2966 ), .C(\U1/aes_core/SB2/n2965 ), .D(
        \U1/aes_core/SB2/n3245 ), .Y(\U1/aes_core/SB2/n2974 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U152  ( .A0(\U1/aes_core/SB2/n2968 ), 
        .A1(\U1/aes_core/SB2/n3212 ), .B0(\U1/aes_core/SB2/n3130 ), .Y(
        \U1/aes_core/SB2/n2970 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U149  ( .A(\U1/aes_core/SB2/n3186 ), .B(
        \U1/aes_core/SB2/n3233 ), .Y(\U1/aes_core/SB2/n3197 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U148  ( .A0(\U1/aes_core/SB2/n3076 ), 
        .A1(\U1/aes_core/SB2/n3255 ), .B0(\U1/aes_core/SB2/n3197 ), .B1(
        \U1/aes_core/SB2/n3208 ), .C0(\U1/aes_core/SB2/n3249 ), .C1(
        \U1/aes_core/SB2/n3258 ), .Y(\U1/aes_core/SB2/n2972 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U147  ( .A(\U1/aes_core/SB2/n2977 ), .B(
        \U1/aes_core/SB2/n2976 ), .C(\U1/aes_core/SB2/n2975 ), .D(
        \U1/aes_core/SB2/n2974 ), .E(\U1/aes_core/SB2/n2973 ), .F(
        \U1/aes_core/SB2/n2972 ), .Y(\U1/aes_core/SB2/n3160 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U146  ( .AN(\U1/aes_core/SB2/n2981 ), 
        .B(\U1/aes_core/SB2/n2980 ), .C(\U1/aes_core/SB2/n2979 ), .D(
        \U1/aes_core/SB2/n2978 ), .Y(\U1/aes_core/SB2/n2991 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB2/U145  ( .A0(\U1/aes_core/SB2/n3243 ), 
        .A1(\U1/aes_core/SB2/n3153 ), .B0(\U1/aes_core/SB2/n3238 ), .B1(
        \U1/aes_core/SB2/n3152 ), .C0(\U1/aes_core/SB2/n2982 ), .C1(
        \U1/aes_core/SB2/n3253 ), .Y(\U1/aes_core/SB2/n2990 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U144  ( .A0(\U1/aes_core/SB2/n3207 ), 
        .A1(\U1/aes_core/SB2/n3113 ), .B0(\U1/aes_core/SB2/n2983 ), .B1(
        \U1/aes_core/SB2/n3076 ), .Y(\U1/aes_core/SB2/n2984 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U143  ( .A0(\U1/aes_core/SB2/n3130 ), 
        .A1(\U1/aes_core/SB2/n3147 ), .B0(\U1/aes_core/SB2/n3146 ), .B1(
        \U1/aes_core/SB2/n3210 ), .C0(\U1/aes_core/SB2/n2984 ), .Y(
        \U1/aes_core/SB2/n2989 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U142  ( .A(\U1/aes_core/SB2/n3218 ), .B(
        \U1/aes_core/SB2/n3257 ), .Y(\U1/aes_core/SB2/n2986 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U141  ( .A0(\U1/aes_core/SB2/n3068 ), 
        .A1(\U1/aes_core/SB2/n2987 ), .B0(\U1/aes_core/SB2/n3239 ), .B1(
        \U1/aes_core/SB2/n2986 ), .C0(\U1/aes_core/SB2/n2985 ), .Y(
        \U1/aes_core/SB2/n2988 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U140  ( .AN(\U1/aes_core/SB2/n2991 ), 
        .B(\U1/aes_core/SB2/n2990 ), .C(\U1/aes_core/SB2/n2989 ), .D(
        \U1/aes_core/SB2/n2988 ), .Y(\U1/aes_core/SB2/n3205 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U139  ( .A(\U1/aes_core/SB2/n2992 ), .Y(
        \U1/aes_core/SB2/n3008 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U138  ( .A0(\U1/aes_core/SB2/n3097 ), 
        .A1(\U1/aes_core/SB2/n3166 ), .B0(\U1/aes_core/SB2/n2993 ), .Y(
        \U1/aes_core/SB2/n3007 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U137  ( .A0(\U1/aes_core/SB2/n3239 ), 
        .A1(\U1/aes_core/SB2/n3238 ), .B0(\U1/aes_core/SB2/n3209 ), .B1(
        \U1/aes_core/SB2/n2994 ), .Y(\U1/aes_core/SB2/n2995 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U136  ( .A0(\U1/aes_core/SB2/n3220 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3236 ), .B1(
        \U1/aes_core/SB2/n3248 ), .C0(\U1/aes_core/SB2/n2995 ), .Y(
        \U1/aes_core/SB2/n3006 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U135  ( .A(\U1/aes_core/SB2/n2999 ), .B(
        \U1/aes_core/SB2/n2998 ), .C(\U1/aes_core/SB2/n2997 ), .D(
        \U1/aes_core/SB2/n2996 ), .Y(\U1/aes_core/SB2/n3005 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U134  ( .AN(\U1/aes_core/SB2/n3003 ), 
        .B(\U1/aes_core/SB2/n3002 ), .C(\U1/aes_core/SB2/n3001 ), .D(
        \U1/aes_core/SB2/n3000 ), .Y(\U1/aes_core/SB2/n3004 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U133  ( .A(\U1/aes_core/SB2/n3009 ), .B(
        \U1/aes_core/SB2/n3008 ), .C(\U1/aes_core/SB2/n3007 ), .D(
        \U1/aes_core/SB2/n3006 ), .E(\U1/aes_core/SB2/n3005 ), .F(
        \U1/aes_core/SB2/n3004 ), .Y(\U1/aes_core/SB2/n3109 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U132  ( .A0(\U1/aes_core/SB2/n3196 ), 
        .A1(\U1/aes_core/SB2/n3113 ), .B0(\U1/aes_core/SB2/n3010 ), .Y(
        \U1/aes_core/SB2/n3025 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U131  ( .AN(\U1/aes_core/SB2/n3014 ), 
        .B(\U1/aes_core/SB2/n3013 ), .C(\U1/aes_core/SB2/n3012 ), .D(
        \U1/aes_core/SB2/n3011 ), .Y(\U1/aes_core/SB2/n3024 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U130  ( .A(\U1/aes_core/SB2/n3230 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3244 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U129  ( .A(\U1/aes_core/SB2/n3017 ), .B(
        \U1/aes_core/SB2/n3016 ), .C(\U1/aes_core/SB2/n3015 ), .D(
        \U1/aes_core/SB2/n3244 ), .Y(\U1/aes_core/SB2/n3023 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U128  ( .A(\U1/aes_core/SB2/n3021 ), .B(
        \U1/aes_core/SB2/n3020 ), .C(\U1/aes_core/SB2/n3019 ), .D(
        \U1/aes_core/SB2/n3018 ), .Y(\U1/aes_core/SB2/n3022 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U127  ( .A(\U1/aes_core/SB2/n3027 ), .B(
        \U1/aes_core/SB2/n3026 ), .C(\U1/aes_core/SB2/n3025 ), .D(
        \U1/aes_core/SB2/n3024 ), .E(\U1/aes_core/SB2/n3023 ), .F(
        \U1/aes_core/SB2/n3022 ), .Y(\U1/aes_core/SB2/n3133 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U126  ( .AN(\U1/aes_core/SB2/n3031 ), 
        .B(\U1/aes_core/SB2/n3030 ), .C(\U1/aes_core/SB2/n3029 ), .D(
        \U1/aes_core/SB2/n3028 ), .Y(\U1/aes_core/SB2/n3040 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U125  ( .A(\U1/aes_core/SB2/n3035 ), .B(
        \U1/aes_core/SB2/n3034 ), .C(\U1/aes_core/SB2/n3033 ), .D(
        \U1/aes_core/SB2/n3032 ), .Y(\U1/aes_core/SB2/n3039 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U124  ( .A(\U1/aes_core/SB2/n3195 ), .B(
        \U1/aes_core/SB2/n3231 ), .C(\U1/aes_core/SB2/n3233 ), .Y(
        \U1/aes_core/SB2/n3037 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U123  ( .A0(\U1/aes_core/SB2/n3037 ), 
        .A1(\U1/aes_core/SB2/n3221 ), .B0(\U1/aes_core/SB2/n3076 ), .B1(
        \U1/aes_core/SB2/n3257 ), .C0(\U1/aes_core/SB2/n3036 ), .Y(
        \U1/aes_core/SB2/n3038 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U122  ( .A(\U1/aes_core/SB2/n3043 ), .B(
        \U1/aes_core/SB2/n3042 ), .C(\U1/aes_core/SB2/n3041 ), .D(
        \U1/aes_core/SB2/n3040 ), .E(\U1/aes_core/SB2/n3039 ), .F(
        \U1/aes_core/SB2/n3038 ), .Y(\U1/aes_core/SB2/n3181 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U121  ( .A0(\U1/aes_core/SB2/n3076 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3044 ), .Y(
        \U1/aes_core/SB2/n3058 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U120  ( .A0(\U1/aes_core/SB2/n3185 ), 
        .A1(\U1/aes_core/SB2/n3187 ), .B0(\U1/aes_core/SB2/n3242 ), .B1(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3045 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U119  ( .A0(\U1/aes_core/SB2/n3096 ), 
        .A1(\U1/aes_core/SB2/n3184 ), .B0(\U1/aes_core/SB2/n3097 ), .B1(
        \U1/aes_core/SB2/n3161 ), .C0(\U1/aes_core/SB2/n3045 ), .Y(
        \U1/aes_core/SB2/n3057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U118  ( .A(\U1/aes_core/SB2/n3046 ), .Y(
        \U1/aes_core/SB2/n3049 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U117  ( .AN(\U1/aes_core/SB2/n3050 ), 
        .B(\U1/aes_core/SB2/n3049 ), .C(\U1/aes_core/SB2/n3048 ), .D(
        \U1/aes_core/SB2/n3047 ), .Y(\U1/aes_core/SB2/n3056 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U116  ( .A(\U1/aes_core/SB2/n3054 ), .B(
        \U1/aes_core/SB2/n3053 ), .C(\U1/aes_core/SB2/n3052 ), .D(
        \U1/aes_core/SB2/n3051 ), .Y(\U1/aes_core/SB2/n3055 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U115  ( .A(\U1/aes_core/SB2/n3060 ), .B(
        \U1/aes_core/SB2/n3059 ), .C(\U1/aes_core/SB2/n3058 ), .D(
        \U1/aes_core/SB2/n3057 ), .E(\U1/aes_core/SB2/n3056 ), .F(
        \U1/aes_core/SB2/n3055 ), .Y(\U1/aes_core/SB2/n3140 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U114  ( .A0(\U1/aes_core/SB2/n3231 ), 
        .A1(\U1/aes_core/SB2/n3061 ), .B0(\U1/aes_core/SB2/n3241 ), .B1(
        \U1/aes_core/SB2/n3187 ), .Y(\U1/aes_core/SB2/n3062 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U113  ( .A0(\U1/aes_core/SB2/n3113 ), 
        .A1(\U1/aes_core/SB2/n3258 ), .B0(\U1/aes_core/SB2/n3063 ), .B1(
        \U1/aes_core/SB2/n3248 ), .C0(\U1/aes_core/SB2/n3062 ), .Y(
        \U1/aes_core/SB2/n3075 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U112  ( .AN(\U1/aes_core/SB2/n3067 ), 
        .B(\U1/aes_core/SB2/n3066 ), .C(\U1/aes_core/SB2/n3065 ), .D(
        \U1/aes_core/SB2/n3064 ), .Y(\U1/aes_core/SB2/n3074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U111  ( .A0(\U1/aes_core/SB2/n3251 ), 
        .A1(\U1/aes_core/SB2/n3068 ), .B0(\U1/aes_core/SB2/n3242 ), .Y(
        \U1/aes_core/SB2/n3072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U110  ( .A(\U1/aes_core/SB2/n3218 ), .B(
        \U1/aes_core/SB2/n3223 ), .Y(\U1/aes_core/SB2/n3069 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U109  ( .A0(\U1/aes_core/SB2/n3194 ), 
        .A1(\U1/aes_core/SB2/n3069 ), .B0(\U1/aes_core/SB2/n3195 ), .B1(
        \U1/aes_core/SB2/n3141 ), .Y(\U1/aes_core/SB2/n3070 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U108  ( .A(\U1/aes_core/SB2/n3072 ), .B(
        \U1/aes_core/SB2/n3071 ), .C(\U1/aes_core/SB2/n3070 ), .Y(
        \U1/aes_core/SB2/n3073 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U107  ( .A(\U1/aes_core/SB2/n3133 ), .B(
        \U1/aes_core/SB2/n3181 ), .C(\U1/aes_core/SB2/n3140 ), .D(
        \U1/aes_core/SB2/n3075 ), .E(\U1/aes_core/SB2/n3074 ), .F(
        \U1/aes_core/SB2/n3073 ), .Y(\U1/aes_core/SB2/n3227 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U106  ( .A(\U1/aes_core/SB2/n3160 ), .B(
        \U1/aes_core/SB2/n3205 ), .C(\U1/aes_core/SB2/n3109 ), .D(
        \U1/aes_core/SB2/n3227 ), .Y(\U1/aes_core/SB2/n3089 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U105  ( .A0(\U1/aes_core/SB2/n3207 ), 
        .A1(\U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3076 ), .B1(
        \U1/aes_core/SB2/n3223 ), .Y(\U1/aes_core/SB2/n3077 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U104  ( .A0(\U1/aes_core/SB2/n3212 ), 
        .A1(\U1/aes_core/SB2/n3230 ), .B0(\U1/aes_core/SB2/n3243 ), .B1(
        \U1/aes_core/SB2/n3251 ), .C0(\U1/aes_core/SB2/n3077 ), .Y(
        \U1/aes_core/SB2/n3088 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U103  ( .A(\U1/aes_core/SB2/n3078 ), .Y(
        \U1/aes_core/SB2/n3081 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U102  ( .A0(\U1/aes_core/SB2/n3079 ), 
        .A1(\U1/aes_core/SB2/n3184 ), .B0(\U1/aes_core/SB2/n3112 ), .B1(
        \U1/aes_core/SB2/n3164 ), .Y(\U1/aes_core/SB2/n3080 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U101  ( .A0(\U1/aes_core/SB2/n3231 ), 
        .A1(\U1/aes_core/SB2/n3081 ), .B0(\U1/aes_core/SB2/n3213 ), .B1(
        \U1/aes_core/SB2/n3162 ), .C0(\U1/aes_core/SB2/n3080 ), .Y(
        \U1/aes_core/SB2/n3087 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U100  ( .A0(\U1/aes_core/SB2/n3253 ), 
        .A1(\U1/aes_core/SB2/n3130 ), .B0(\U1/aes_core/SB2/n3233 ), .Y(
        \U1/aes_core/SB2/n3085 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB2/U99  ( .A(\U1/aes_core/SB2/n3085 ), .B(
        \U1/aes_core/SB2/n3084 ), .C(\U1/aes_core/SB2/n3083 ), .D(
        \U1/aes_core/SB2/n3082 ), .Y(\U1/aes_core/SB2/n3086 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U98  ( .AN(\U1/aes_core/SB2/n3089 ), .B(
        \U1/aes_core/SB2/n3088 ), .C(\U1/aes_core/SB2/n3087 ), .D(
        \U1/aes_core/SB2/n3086 ), .Y(\U1/aes_core/sb2 [3]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U97  ( .A0(\U1/aes_core/SB2/n3104 ), .A1(
        \U1/aes_core/SB2/n3219 ), .B0(\U1/aes_core/SB2/n3163 ), .Y(
        \U1/aes_core/SB2/n3101 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U96  ( .A(\U1/aes_core/SB2/n3092 ), .B(
        \U1/aes_core/SB2/n3091 ), .C(\U1/aes_core/SB2/n3090 ), .Y(
        \U1/aes_core/SB2/n3100 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U95  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3242 ), .Y(\U1/aes_core/SB2/n3095 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U94  ( .A(\U1/aes_core/SB2/n3213 ), .B(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3093 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U93  ( .A0(\U1/aes_core/SB2/n3095 ), 
        .A1(\U1/aes_core/SB2/n3094 ), .B0(\U1/aes_core/SB2/n3093 ), .B1(
        \U1/aes_core/SB2/n3236 ), .C0(\U1/aes_core/SB2/n3219 ), .C1(
        \U1/aes_core/SB2/n3145 ), .Y(\U1/aes_core/SB2/n3099 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U92  ( .A0(\U1/aes_core/SB2/n3196 ), 
        .A1(\U1/aes_core/SB2/n3097 ), .B0(\U1/aes_core/SB2/n3258 ), .B1(
        \U1/aes_core/SB2/n3248 ), .C0(\U1/aes_core/SB2/n3221 ), .C1(
        \U1/aes_core/SB2/n3096 ), .Y(\U1/aes_core/SB2/n3098 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U91  ( .A(\U1/aes_core/SB2/n3103 ), .B(
        \U1/aes_core/SB2/n3102 ), .C(\U1/aes_core/SB2/n3101 ), .D(
        \U1/aes_core/SB2/n3100 ), .E(\U1/aes_core/SB2/n3099 ), .F(
        \U1/aes_core/SB2/n3098 ), .Y(\U1/aes_core/SB2/n3228 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB2/U90  ( .A0(\U1/aes_core/SB2/n3104 ), .A1(
        \U1/aes_core/SB2/n3113 ), .B0(\U1/aes_core/SB2/n3184 ), .Y(
        \U1/aes_core/SB2/n3139 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB2/U89  ( .A0(\U1/aes_core/SB2/n3208 ), .A1(
        \U1/aes_core/SB2/n3221 ), .A2(\U1/aes_core/SB2/n3161 ), .B0(
        \U1/aes_core/SB2/n3237 ), .Y(\U1/aes_core/SB2/n3138 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U88  ( .A(\U1/aes_core/SB2/n3108 ), .B(
        \U1/aes_core/SB2/n3107 ), .C(\U1/aes_core/SB2/n3106 ), .D(
        \U1/aes_core/SB2/n3105 ), .Y(\U1/aes_core/SB2/n3135 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U87  ( .A(\U1/aes_core/SB2/n3109 ), .Y(
        \U1/aes_core/SB2/n3132 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U86  ( .A(\U1/aes_core/SB2/n3110 ), .Y(
        \U1/aes_core/SB2/n3126 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB2/U85  ( .A0(\U1/aes_core/SB2/n3112 ), 
        .A1(\U1/aes_core/SB2/n3249 ), .B0N(\U1/aes_core/SB2/n3111 ), .Y(
        \U1/aes_core/SB2/n3125 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U84  ( .A0(\U1/aes_core/SB2/n3256 ), 
        .A1(\U1/aes_core/SB2/n3113 ), .B0(\U1/aes_core/SB2/n3163 ), .B1(
        \U1/aes_core/SB2/n3223 ), .C0(\U1/aes_core/SB2/n3237 ), .C1(
        \U1/aes_core/SB2/n3258 ), .Y(\U1/aes_core/SB2/n3124 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U83  ( .AN(\U1/aes_core/SB2/n3117 ), .B(
        \U1/aes_core/SB2/n3116 ), .C(\U1/aes_core/SB2/n3115 ), .D(
        \U1/aes_core/SB2/n3114 ), .Y(\U1/aes_core/SB2/n3123 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U82  ( .A(\U1/aes_core/SB2/n3121 ), .B(
        \U1/aes_core/SB2/n3120 ), .C(\U1/aes_core/SB2/n3119 ), .D(
        \U1/aes_core/SB2/n3118 ), .Y(\U1/aes_core/SB2/n3122 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U81  ( .A(\U1/aes_core/SB2/n3127 ), .B(
        \U1/aes_core/SB2/n3126 ), .C(\U1/aes_core/SB2/n3125 ), .D(
        \U1/aes_core/SB2/n3124 ), .E(\U1/aes_core/SB2/n3123 ), .F(
        \U1/aes_core/SB2/n3122 ), .Y(\U1/aes_core/SB2/n3128 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U80  ( .A(\U1/aes_core/SB2/n3128 ), .Y(
        \U1/aes_core/SB2/n3206 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U79  ( .A0(\U1/aes_core/SB2/n3196 ), .A1(
        \U1/aes_core/SB2/n3218 ), .B0(\U1/aes_core/SB2/n3258 ), .B1(
        \U1/aes_core/SB2/n3257 ), .Y(\U1/aes_core/SB2/n3129 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U78  ( .A0(\U1/aes_core/SB2/n3186 ), 
        .A1(\U1/aes_core/SB2/n3130 ), .B0(\U1/aes_core/SB2/n3210 ), .B1(
        \U1/aes_core/SB2/n3232 ), .C0(\U1/aes_core/SB2/n3129 ), .Y(
        \U1/aes_core/SB2/n3131 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U77  ( .AN(\U1/aes_core/SB2/n3133 ), .B(
        \U1/aes_core/SB2/n3132 ), .C(\U1/aes_core/SB2/n3206 ), .D(
        \U1/aes_core/SB2/n3131 ), .Y(\U1/aes_core/SB2/n3134 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U76  ( .A(\U1/aes_core/SB2/n3139 ), .B(
        \U1/aes_core/SB2/n3138 ), .C(\U1/aes_core/SB2/n3137 ), .D(
        \U1/aes_core/SB2/n3136 ), .E(\U1/aes_core/SB2/n3135 ), .F(
        \U1/aes_core/SB2/n3134 ), .Y(\U1/aes_core/SB2/n3204 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U75  ( .A(\U1/aes_core/SB2/n3140 ), .Y(
        \U1/aes_core/SB2/n3144 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U74  ( .A0(\U1/aes_core/SB2/n3142 ), .A1(
        \U1/aes_core/SB2/n3141 ), .B0(\U1/aes_core/SB2/n3188 ), .B1(
        \U1/aes_core/SB2/n3147 ), .Y(\U1/aes_core/SB2/n3143 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U73  ( .A0(\U1/aes_core/SB2/n3237 ), 
        .A1(\U1/aes_core/SB2/n3145 ), .B0(\U1/aes_core/SB2/n3144 ), .C0(
        \U1/aes_core/SB2/n3143 ), .Y(\U1/aes_core/SB2/n3159 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U72  ( .A0(\U1/aes_core/SB2/n3146 ), .A1(
        \U1/aes_core/SB2/n3209 ), .B0(\U1/aes_core/SB2/n3238 ), .Y(
        \U1/aes_core/SB2/n3151 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U71  ( .A0(\U1/aes_core/SB2/n3147 ), .A1(
        \U1/aes_core/SB2/n3212 ), .B0(\U1/aes_core/SB2/n3241 ), .Y(
        \U1/aes_core/SB2/n3150 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U70  ( .A(\U1/aes_core/SB2/n3151 ), .B(
        \U1/aes_core/SB2/n3150 ), .C(\U1/aes_core/SB2/n3149 ), .D(
        \U1/aes_core/SB2/n3148 ), .Y(\U1/aes_core/SB2/n3158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U69  ( .A(\U1/aes_core/SB2/n3189 ), .B(
        \U1/aes_core/SB2/n3152 ), .Y(\U1/aes_core/SB2/n3156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U68  ( .A(\U1/aes_core/SB2/n3153 ), .B(
        \U1/aes_core/SB2/n3194 ), .Y(\U1/aes_core/SB2/n3155 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U67  ( .A0(\U1/aes_core/SB2/n3156 ), 
        .A1(\U1/aes_core/SB2/n3255 ), .B0(\U1/aes_core/SB2/n3155 ), .B1(
        \U1/aes_core/SB2/n3219 ), .C0(\U1/aes_core/SB2/n3154 ), .C1(
        \U1/aes_core/SB2/n3220 ), .Y(\U1/aes_core/SB2/n3157 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U66  ( .A(\U1/aes_core/SB2/n3228 ), .B(
        \U1/aes_core/SB2/n3204 ), .C(\U1/aes_core/SB2/n3160 ), .D(
        \U1/aes_core/SB2/n3159 ), .E(\U1/aes_core/SB2/n3158 ), .F(
        \U1/aes_core/SB2/n3157 ), .Y(\U1/aes_core/sb2 [4]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U65  ( .A1N(\U1/aes_core/SB2/n3162 ), 
        .A0(\U1/aes_core/SB2/n3161 ), .B0(\U1/aes_core/SB2/n3218 ), .Y(
        \U1/aes_core/SB2/n3178 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U64  ( .A(\U1/aes_core/SB2/n3231 ), .B(
        \U1/aes_core/SB2/n3212 ), .Y(\U1/aes_core/SB2/n3165 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U63  ( .A0(\U1/aes_core/SB2/n3255 ), 
        .A1(\U1/aes_core/SB2/n3166 ), .B0(\U1/aes_core/SB2/n3165 ), .B1(
        \U1/aes_core/SB2/n3258 ), .C0(\U1/aes_core/SB2/n3164 ), .C1(
        \U1/aes_core/SB2/n3163 ), .Y(\U1/aes_core/SB2/n3177 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U62  ( .A(\U1/aes_core/SB2/n3167 ), .Y(
        \U1/aes_core/SB2/n3170 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U61  ( .AN(\U1/aes_core/SB2/n3171 ), .B(
        \U1/aes_core/SB2/n3170 ), .C(\U1/aes_core/SB2/n3169 ), .D(
        \U1/aes_core/SB2/n3168 ), .Y(\U1/aes_core/SB2/n3176 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U60  ( .A(\U1/aes_core/SB2/n3174 ), .B(
        \U1/aes_core/SB2/n3173 ), .C(\U1/aes_core/SB2/n3172 ), .Y(
        \U1/aes_core/SB2/n3175 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U59  ( .A(\U1/aes_core/SB2/n3180 ), .B(
        \U1/aes_core/SB2/n3179 ), .C(\U1/aes_core/SB2/n3178 ), .D(
        \U1/aes_core/SB2/n3177 ), .E(\U1/aes_core/SB2/n3176 ), .F(
        \U1/aes_core/SB2/n3175 ), .Y(\U1/aes_core/SB2/n3229 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U58  ( .A(\U1/aes_core/SB2/n3181 ), .Y(
        \U1/aes_core/SB2/n3183 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U57  ( .A0(\U1/aes_core/SB2/n3242 ), .A1(
        \U1/aes_core/SB2/n3239 ), .B0(\U1/aes_core/SB2/n3243 ), .B1(
        \U1/aes_core/SB2/n3241 ), .Y(\U1/aes_core/SB2/n3182 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U56  ( .A0(\U1/aes_core/SB2/n3218 ), 
        .A1(\U1/aes_core/SB2/n3184 ), .B0(\U1/aes_core/SB2/n3183 ), .C0(
        \U1/aes_core/SB2/n3182 ), .Y(\U1/aes_core/SB2/n3203 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U55  ( .A0(\U1/aes_core/SB2/n3186 ), .A1(
        \U1/aes_core/SB2/n3242 ), .B0(\U1/aes_core/SB2/n3185 ), .Y(
        \U1/aes_core/SB2/n3192 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U54  ( .A0(\U1/aes_core/SB2/n3189 ), .A1(
        \U1/aes_core/SB2/n3188 ), .B0(\U1/aes_core/SB2/n3187 ), .Y(
        \U1/aes_core/SB2/n3191 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U53  ( .AN(\U1/aes_core/SB2/n3193 ), .B(
        \U1/aes_core/SB2/n3192 ), .C(\U1/aes_core/SB2/n3191 ), .D(
        \U1/aes_core/SB2/n3190 ), .Y(\U1/aes_core/SB2/n3202 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U52  ( .A0(\U1/aes_core/SB2/n3238 ), .A1(
        \U1/aes_core/SB2/n3195 ), .B0(\U1/aes_core/SB2/n3194 ), .Y(
        \U1/aes_core/SB2/n3199 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB2/U51  ( .A0(\U1/aes_core/SB2/n3220 ), .A1(
        \U1/aes_core/SB2/n3197 ), .B0(\U1/aes_core/SB2/n3257 ), .B1(
        \U1/aes_core/SB2/n3196 ), .Y(\U1/aes_core/SB2/n3198 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U50  ( .A0(\U1/aes_core/SB2/n3200 ), 
        .A1(\U1/aes_core/SB2/n3219 ), .B0(\U1/aes_core/SB2/n3199 ), .C0(
        \U1/aes_core/SB2/n3198 ), .Y(\U1/aes_core/SB2/n3201 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U49  ( .A(\U1/aes_core/SB2/n3229 ), .B(
        \U1/aes_core/SB2/n3205 ), .C(\U1/aes_core/SB2/n3204 ), .D(
        \U1/aes_core/SB2/n3203 ), .E(\U1/aes_core/SB2/n3202 ), .F(
        \U1/aes_core/SB2/n3201 ), .Y(\U1/aes_core/sb2 [5]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U48  ( .A0(\U1/aes_core/SB2/n3208 ), 
        .A1(\U1/aes_core/SB2/n3248 ), .B0(\U1/aes_core/SB2/n3207 ), .B1(
        \U1/aes_core/SB2/n3255 ), .C0(\U1/aes_core/SB2/n3206 ), .Y(
        \U1/aes_core/SB2/n3226 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U47  ( .A0(\U1/aes_core/SB2/n3209 ), .A1(
        \U1/aes_core/SB2/n3253 ), .B0(\U1/aes_core/SB2/n3242 ), .Y(
        \U1/aes_core/SB2/n3217 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U46  ( .A0(\U1/aes_core/SB2/n3233 ), .A1(
        \U1/aes_core/SB2/n3210 ), .B0(\U1/aes_core/SB2/n3241 ), .Y(
        \U1/aes_core/SB2/n3216 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U45  ( .A0(\U1/aes_core/SB2/n3213 ), .A1(
        \U1/aes_core/SB2/n3212 ), .B0(\U1/aes_core/SB2/n3211 ), .Y(
        \U1/aes_core/SB2/n3215 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U44  ( .A(\U1/aes_core/SB2/n3217 ), .B(
        \U1/aes_core/SB2/n3216 ), .C(\U1/aes_core/SB2/n3215 ), .D(
        \U1/aes_core/SB2/n3214 ), .Y(\U1/aes_core/SB2/n3225 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U43  ( .A(\U1/aes_core/SB2/n3248 ), .B(
        \U1/aes_core/SB2/n3218 ), .Y(\U1/aes_core/SB2/n3250 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB2/U42  ( .A(\U1/aes_core/SB2/n3238 ), .B(
        \U1/aes_core/SB2/n3250 ), .Y(\U1/aes_core/SB2/n3222 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U41  ( .A0(\U1/aes_core/SB2/n3236 ), 
        .A1(\U1/aes_core/SB2/n3223 ), .B0(\U1/aes_core/SB2/n3222 ), .B1(
        \U1/aes_core/SB2/n3221 ), .C0(\U1/aes_core/SB2/n3220 ), .C1(
        \U1/aes_core/SB2/n3219 ), .Y(\U1/aes_core/SB2/n3224 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U40  ( .A(\U1/aes_core/SB2/n3229 ), .B(
        \U1/aes_core/SB2/n3228 ), .C(\U1/aes_core/SB2/n3227 ), .D(
        \U1/aes_core/SB2/n3226 ), .E(\U1/aes_core/SB2/n3225 ), .F(
        \U1/aes_core/SB2/n3224 ), .Y(\U1/aes_core/sb2 [6]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U39  ( .A0(\U1/aes_core/SB2/n3233 ), .A1(
        \U1/aes_core/SB2/n3232 ), .B0(\U1/aes_core/SB2/n3231 ), .B1(
        \U1/aes_core/SB2/n3230 ), .Y(\U1/aes_core/SB2/n3234 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB2/U38  ( .A0(\U1/aes_core/SB2/n3237 ), 
        .A1(\U1/aes_core/SB2/n3236 ), .B0(\U1/aes_core/SB2/n3235 ), .C0(
        \U1/aes_core/SB2/n3234 ), .Y(\U1/aes_core/SB2/n3261 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB2/U37  ( .A1N(\U1/aes_core/SB2/n3240 ), 
        .A0(\U1/aes_core/SB2/n3239 ), .B0(\U1/aes_core/SB2/n3238 ), .Y(
        \U1/aes_core/SB2/n3247 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U36  ( .A0(\U1/aes_core/SB2/n3243 ), .A1(
        \U1/aes_core/SB2/n3242 ), .B0(\U1/aes_core/SB2/n3241 ), .Y(
        \U1/aes_core/SB2/n3246 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U35  ( .A(\U1/aes_core/SB2/n3247 ), .B(
        \U1/aes_core/SB2/n3246 ), .C(\U1/aes_core/SB2/n3245 ), .D(
        \U1/aes_core/SB2/n3244 ), .Y(\U1/aes_core/SB2/n3260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U34  ( .A(\U1/aes_core/SB2/n3249 ), .B(
        \U1/aes_core/SB2/n3248 ), .Y(\U1/aes_core/SB2/n3252 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U33  ( .A0(\U1/aes_core/SB2/n3253 ), .A1(
        \U1/aes_core/SB2/n3252 ), .B0(\U1/aes_core/SB2/n3251 ), .B1(
        \U1/aes_core/SB2/n3250 ), .Y(\U1/aes_core/SB2/n3254 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U32  ( .A0(\U1/aes_core/SB2/n3258 ), 
        .A1(\U1/aes_core/SB2/n3257 ), .B0(\U1/aes_core/SB2/n3256 ), .B1(
        \U1/aes_core/SB2/n3255 ), .C0(\U1/aes_core/SB2/n3254 ), .Y(
        \U1/aes_core/SB2/n3259 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U31  ( .A(\U1/aes_core/SB2/n3264 ), .B(
        \U1/aes_core/SB2/n3263 ), .C(\U1/aes_core/SB2/n3262 ), .D(
        \U1/aes_core/SB2/n3261 ), .E(\U1/aes_core/SB2/n3260 ), .F(
        \U1/aes_core/SB2/n3259 ), .Y(\U1/aes_core/sb2 [7]) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U30  ( .A(\U1/aes_core/SB2/n3267 ), .B(
        \U1/aes_core/SB2/n3266 ), .C(\U1/aes_core/SB2/n3265 ), .Y(
        \U1/aes_core/SB2/n3290 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U29  ( .A0(\U1/aes_core/SB2/n3268 ), .A1(
        \U1/aes_core/SB2/n3324 ), .B0(\U1/aes_core/SB2/n3340 ), .Y(
        \U1/aes_core/SB2/n3273 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U28  ( .A0(\U1/aes_core/SB2/n3333 ), .A1(
        \U1/aes_core/SB2/n3270 ), .B0(\U1/aes_core/SB2/n3269 ), .B1(
        \U1/aes_core/SB2/n3334 ), .Y(\U1/aes_core/SB2/n3271 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U27  ( .A(\U1/aes_core/SB2/n3273 ), .B(
        \U1/aes_core/SB2/n3272 ), .C(\U1/aes_core/SB2/n3271 ), .Y(
        \U1/aes_core/SB2/n3289 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB2/U26  ( .A0(\U1/aes_core/SB2/n3276 ), .A1(
        \U1/aes_core/SB2/n3299 ), .B0(\U1/aes_core/SB2/n3275 ), .B1(
        \U1/aes_core/SB2/n3274 ), .Y(\U1/aes_core/SB2/n3277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB2/U25  ( .A0(\U1/aes_core/SB2/n3281 ), 
        .A1(\U1/aes_core/SB2/n3280 ), .B0(\U1/aes_core/SB2/n3279 ), .B1(
        \U1/aes_core/SB2/n3278 ), .C0(\U1/aes_core/SB2/n3277 ), .Y(
        \U1/aes_core/SB2/n3288 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U24  ( .A(\U1/aes_core/SB2/n3329 ), .B(
        \U1/aes_core/SB2/n3282 ), .Y(\U1/aes_core/SB2/n3283 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U23  ( .AN(\U1/aes_core/SB2/n3286 ), .B(
        \U1/aes_core/SB2/n3285 ), .C(\U1/aes_core/SB2/n3284 ), .D(
        \U1/aes_core/SB2/n3283 ), .Y(\U1/aes_core/SB2/n3287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U22  ( .A(\U1/aes_core/SB2/n3292 ), .B(
        \U1/aes_core/SB2/n3291 ), .C(\U1/aes_core/SB2/n3290 ), .D(
        \U1/aes_core/SB2/n3289 ), .E(\U1/aes_core/SB2/n3288 ), .F(
        \U1/aes_core/SB2/n3287 ), .Y(\U1/aes_core/SB2/n3351 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB2/U21  ( .A(\U1/aes_core/SB2/n3295 ), .B(
        \U1/aes_core/SB2/n3294 ), .C(\U1/aes_core/SB2/n3293 ), .D(
        \U1/aes_core/SB2/n3351 ), .Y(\U1/aes_core/SB2/n3320 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U20  ( .A0(\U1/aes_core/SB2/n3297 ), .A1(
        \U1/aes_core/SB2/n3308 ), .B0(\U1/aes_core/SB2/n3344 ), .B1(
        \U1/aes_core/SB2/n3296 ), .Y(\U1/aes_core/SB2/n3298 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U19  ( .A0(\U1/aes_core/SB2/n3322 ), 
        .A1(\U1/aes_core/SB2/n3334 ), .B0(\U1/aes_core/SB2/n3325 ), .B1(
        \U1/aes_core/SB2/n3299 ), .C0(\U1/aes_core/SB2/n3298 ), .Y(
        \U1/aes_core/SB2/n3319 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB2/U18  ( .A0(\U1/aes_core/SB2/n3303 ), .A1(
        \U1/aes_core/SB2/n3302 ), .B0(\U1/aes_core/SB2/n3301 ), .B1(
        \U1/aes_core/SB2/n3300 ), .Y(\U1/aes_core/SB2/n3304 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U17  ( .A0(\U1/aes_core/SB2/n3307 ), 
        .A1(\U1/aes_core/SB2/n3306 ), .B0(\U1/aes_core/SB2/n3305 ), .B1(
        \U1/aes_core/SB2/n3330 ), .C0(\U1/aes_core/SB2/n3304 ), .Y(
        \U1/aes_core/SB2/n3318 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB2/U16  ( .A(\U1/aes_core/SB2/n3309 ), .B(
        \U1/aes_core/SB2/n3308 ), .Y(\U1/aes_core/SB2/n3316 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U15  ( .A(\U1/aes_core/SB2/n3310 ), .Y(
        \U1/aes_core/SB2/n3315 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB2/U14  ( .A(\U1/aes_core/SB2/n3313 ), .B(
        \U1/aes_core/SB2/n3312 ), .C(\U1/aes_core/SB2/n3311 ), .Y(
        \U1/aes_core/SB2/n3314 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U13  ( .A0(\U1/aes_core/SB2/n3331 ), 
        .A1(\U1/aes_core/SB2/n3316 ), .B0(\U1/aes_core/SB2/n3323 ), .B1(
        \U1/aes_core/SB2/n3315 ), .C0(\U1/aes_core/SB2/n3314 ), .Y(
        \U1/aes_core/SB2/n3317 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB2/U12  ( .AN(\U1/aes_core/SB2/n3320 ), .B(
        \U1/aes_core/SB2/n3319 ), .C(\U1/aes_core/SB2/n3318 ), .D(
        \U1/aes_core/SB2/n3317 ), .Y(\U1/aes_core/sb2 [8]) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB2/U11  ( .A0(\U1/aes_core/SB2/n3325 ), 
        .A1(\U1/aes_core/SB2/n3324 ), .B0(\U1/aes_core/SB2/n3323 ), .B1(
        \U1/aes_core/SB2/n3322 ), .C0(\U1/aes_core/SB2/n3321 ), .Y(
        \U1/aes_core/SB2/n3326 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB2/U10  ( .A(\U1/aes_core/SB2/n3326 ), .Y(
        \U1/aes_core/SB2/n3350 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U9  ( .A0(\U1/aes_core/SB2/n3339 ), .A1(
        \U1/aes_core/SB2/n3328 ), .B0(\U1/aes_core/SB2/n3327 ), .Y(
        \U1/aes_core/SB2/n3338 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U8  ( .A0(\U1/aes_core/SB2/n3331 ), .A1(
        \U1/aes_core/SB2/n3330 ), .B0(\U1/aes_core/SB2/n3329 ), .Y(
        \U1/aes_core/SB2/n3337 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB2/U7  ( .A0(\U1/aes_core/SB2/n3334 ), .A1(
        \U1/aes_core/SB2/n3333 ), .B0(\U1/aes_core/SB2/n3332 ), .Y(
        \U1/aes_core/SB2/n3336 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB2/U6  ( .A(\U1/aes_core/SB2/n3338 ), .B(
        \U1/aes_core/SB2/n3337 ), .C(\U1/aes_core/SB2/n3336 ), .D(
        \U1/aes_core/SB2/n3335 ), .Y(\U1/aes_core/SB2/n3349 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB2/U5  ( .A(\U1/aes_core/SB2/n3341 ), .B(
        \U1/aes_core/SB2/n3340 ), .C(\U1/aes_core/SB2/n3339 ), .Y(
        \U1/aes_core/SB2/n3345 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB2/U4  ( .A0(\U1/aes_core/SB2/n3347 ), .A1(
        \U1/aes_core/SB2/n3346 ), .B0(\U1/aes_core/SB2/n3345 ), .B1(
        \U1/aes_core/SB2/n3344 ), .C0(\U1/aes_core/SB2/n3343 ), .C1(
        \U1/aes_core/SB2/n3342 ), .Y(\U1/aes_core/SB2/n3348 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB2/U3  ( .A(\U1/aes_core/SB2/n3353 ), .B(
        \U1/aes_core/SB2/n3352 ), .C(\U1/aes_core/SB2/n3351 ), .D(
        \U1/aes_core/SB2/n3350 ), .E(\U1/aes_core/SB2/n3349 ), .F(
        \U1/aes_core/SB2/n3348 ), .Y(\U1/aes_core/sb2 [9]) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U711  ( .A0(\U1/aes_core/SB3/n2971 ), .A1(
        \U1/aes_core/SB3/n3096 ), .B0(\U1/aes_core/SB3/n3094 ), .B1(
        \U1/aes_core/SB3/n3079 ), .C0(\U1/aes_core/SB3/n2970 ), .Y(
        \U1/aes_core/SB3/n2973 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U393  ( .A0(\U1/aes_core/SB3/n2402 ), .A1(
        \U1/aes_core/SB3/n2157 ), .B0(\U1/aes_core/SB3/n2480 ), .B1(
        \U1/aes_core/SB3/n2464 ), .C0(\U1/aes_core/SB3/n2225 ), .Y(
        \U1/aes_core/SB3/n2158 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U391  ( .A0(\U1/aes_core/SB3/n2650 ), .A1(
        \U1/aes_core/SB3/n2775 ), .B0(\U1/aes_core/SB3/n2773 ), .B1(
        \U1/aes_core/SB3/n2758 ), .C0(\U1/aes_core/SB3/n2649 ), .Y(
        \U1/aes_core/SB3/n2652 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U363  ( .A0(\U1/aes_core/SB3/n3145 ), .A1(
        \U1/aes_core/SB3/n2328 ), .B0(\U1/aes_core/SB3/n3223 ), .B1(
        \U1/aes_core/SB3/n3207 ), .C0(\U1/aes_core/SB3/n2993 ), .Y(
        \U1/aes_core/SB3/n2329 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U361  ( .A0(\U1/aes_core/SB3/n2203 ), .A1(
        \U1/aes_core/SB3/n2353 ), .B0(\U1/aes_core/SB3/n2351 ), .B1(
        \U1/aes_core/SB3/n2311 ), .C0(\U1/aes_core/SB3/n2202 ), .Y(
        \U1/aes_core/SB3/n2205 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U301  ( .A0(\U1/aes_core/SB3/n2824 ), .A1(
        \U1/aes_core/SB3/n2604 ), .B0(\U1/aes_core/SB3/n2923 ), .B1(
        \U1/aes_core/SB3/n2907 ), .C0(\U1/aes_core/SB3/n2672 ), .Y(
        \U1/aes_core/SB3/n2605 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U300  ( .A0(\U1/aes_core/SB3/n3145 ), .A1(
        \U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3223 ), .B1(
        \U1/aes_core/SB3/n3221 ), .C0(\U1/aes_core/SB3/n3036 ), .Y(
        \U1/aes_core/SB3/n1742 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U151  ( .A0(\U1/aes_core/SB3/n2402 ), .A1(
        \U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2480 ), .B1(
        \U1/aes_core/SB3/n2478 ), .C0(\U1/aes_core/SB3/n2268 ), .Y(
        \U1/aes_core/SB3/n2144 ) );
  OAI221_X1M_A12TL \U1/aes_core/SB3/U150  ( .A0(\U1/aes_core/SB3/n2824 ), .A1(
        \U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2923 ), .B1(
        \U1/aes_core/SB3/n2921 ), .C0(\U1/aes_core/SB3/n2715 ), .Y(
        \U1/aes_core/SB3/n2591 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1724  ( .A(Dout[7]), .B(Dout[6]), .Y(
        \U1/aes_core/SB3/n1691 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1723  ( .A(Dout[5]), .B(Dout[4]), .Y(
        \U1/aes_core/SB3/n1682 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1722  ( .A(\U1/aes_core/SB3/n1691 ), .B(
        \U1/aes_core/SB3/n1682 ), .Y(\U1/aes_core/SB3/n2328 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1721  ( .A(Dout[1]), .Y(
        \U1/aes_core/SB3/n767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1720  ( .A(Dout[0]), .Y(
        \U1/aes_core/SB3/n385 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1719  ( .A(\U1/aes_core/SB3/n767 ), .B(
        \U1/aes_core/SB3/n385 ), .Y(\U1/aes_core/SB3/n1683 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1718  ( .A(Dout[3]), .B(Dout[2]), .Y(
        \U1/aes_core/SB3/n1703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1717  ( .A(\U1/aes_core/SB3/n1683 ), .B(
        \U1/aes_core/SB3/n1703 ), .Y(\U1/aes_core/SB3/n3207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1716  ( .A(\U1/aes_core/SB3/n2328 ), .B(
        \U1/aes_core/SB3/n3207 ), .Y(\U1/aes_core/SB3/n3014 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U1715  ( .A(Dout[2]), .B(Dout[3]), .Y(
        \U1/aes_core/SB3/n1686 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1714  ( .A(\U1/aes_core/SB3/n1686 ), .B(
        \U1/aes_core/SB3/n1683 ), .Y(\U1/aes_core/SB3/n3145 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1713  ( .A(Dout[7]), .Y(
        \U1/aes_core/SB3/n1203 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1712  ( .A(\U1/aes_core/SB3/n1203 ), .B(
        Dout[6]), .Y(\U1/aes_core/SB3/n1709 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1711  ( .A(\U1/aes_core/SB3/n1709 ), .B(
        \U1/aes_core/SB3/n1682 ), .Y(\U1/aes_core/SB3/n2327 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1710  ( .A(\U1/aes_core/SB3/n3145 ), .B(
        \U1/aes_core/SB3/n2327 ), .Y(\U1/aes_core/SB3/n3111 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1709  ( .A(Dout[3]), .Y(
        \U1/aes_core/SB3/n707 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U1708  ( .A(Dout[2]), .B(
        \U1/aes_core/SB3/n707 ), .Y(\U1/aes_core/SB3/n1684 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1707  ( .A(\U1/aes_core/SB3/n1683 ), .B(
        \U1/aes_core/SB3/n1684 ), .Y(\U1/aes_core/SB3/n3076 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1706  ( .A(\U1/aes_core/SB3/n3076 ), .Y(
        \U1/aes_core/SB3/n3241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1705  ( .A(Dout[4]), .Y(
        \U1/aes_core/SB3/n752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1704  ( .A(\U1/aes_core/SB3/n752 ), .B(
        Dout[5]), .Y(\U1/aes_core/SB3/n1690 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1703  ( .A(Dout[6]), .Y(
        \U1/aes_core/SB3/n1158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1702  ( .A(\U1/aes_core/SB3/n1158 ), .B(
        Dout[7]), .Y(\U1/aes_core/SB3/n1700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1701  ( .A(\U1/aes_core/SB3/n1690 ), .B(
        \U1/aes_core/SB3/n1700 ), .Y(\U1/aes_core/SB3/n3097 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1700  ( .A(\U1/aes_core/SB3/n3097 ), .Y(
        \U1/aes_core/SB3/n3195 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1699  ( .A(\U1/aes_core/SB3/n3241 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n3054 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1698  ( .A(\U1/aes_core/SB3/n2328 ), .Y(
        \U1/aes_core/SB3/n3210 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1697  ( .A(Dout[1]), .B(Dout[0]), .Y(
        \U1/aes_core/SB3/n1687 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1696  ( .A(\U1/aes_core/SB3/n1687 ), .B(
        \U1/aes_core/SB3/n1703 ), .Y(\U1/aes_core/SB3/n3163 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1695  ( .A(\U1/aes_core/SB3/n3163 ), .Y(
        \U1/aes_core/SB3/n3251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1694  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3251 ), .Y(\U1/aes_core/SB3/n3168 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1693  ( .A(\U1/aes_core/SB3/n385 ), .B(
        Dout[1]), .Y(\U1/aes_core/SB3/n1702 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1692  ( .A(\U1/aes_core/SB3/n1684 ), .B(
        \U1/aes_core/SB3/n1702 ), .Y(\U1/aes_core/SB3/n3063 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1691  ( .A(\U1/aes_core/SB3/n3063 ), .Y(
        \U1/aes_core/SB3/n3152 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1690  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3032 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U1689  ( .A(\U1/aes_core/SB3/n3054 ), .B(
        \U1/aes_core/SB3/n3168 ), .C(\U1/aes_core/SB3/n3032 ), .Y(
        \U1/aes_core/SB3/n1722 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1688  ( .A(\U1/aes_core/SB3/n1682 ), .B(
        \U1/aes_core/SB3/n1700 ), .Y(\U1/aes_core/SB3/n3096 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1687  ( .A(\U1/aes_core/SB3/n707 ), .B(
        Dout[2]), .Y(\U1/aes_core/SB3/n1693 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1686  ( .A(\U1/aes_core/SB3/n1693 ), .B(
        \U1/aes_core/SB3/n1702 ), .Y(\U1/aes_core/SB3/n3094 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1685  ( .A(\U1/aes_core/SB3/n3096 ), .B(
        \U1/aes_core/SB3/n3094 ), .Y(\U1/aes_core/SB3/n3009 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1684  ( .A(\U1/aes_core/SB3/n2327 ), .Y(
        \U1/aes_core/SB3/n3212 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1683  ( .A(Dout[5]), .Y(
        \U1/aes_core/SB3/n1030 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1682  ( .A(\U1/aes_core/SB3/n752 ), .B(
        \U1/aes_core/SB3/n1030 ), .Y(\U1/aes_core/SB3/n1701 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1681  ( .A(\U1/aes_core/SB3/n1691 ), .B(
        \U1/aes_core/SB3/n1701 ), .Y(\U1/aes_core/SB3/n3255 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1680  ( .A(\U1/aes_core/SB3/n3255 ), .Y(
        \U1/aes_core/SB3/n3186 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1679  ( .A(\U1/aes_core/SB3/n767 ), .B(
        Dout[0]), .Y(\U1/aes_core/SB3/n1692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1678  ( .A(\U1/aes_core/SB3/n1692 ), .B(
        \U1/aes_core/SB3/n1703 ), .Y(\U1/aes_core/SB3/n3220 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1677  ( .A(\U1/aes_core/SB3/n3220 ), .Y(
        \U1/aes_core/SB3/n3068 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1676  ( .A0(\U1/aes_core/SB3/n3212 ), 
        .A1(\U1/aes_core/SB3/n3186 ), .B0(\U1/aes_core/SB3/n3068 ), .Y(
        \U1/aes_core/SB3/n1621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1675  ( .A(\U1/aes_core/SB3/n1687 ), .B(
        \U1/aes_core/SB3/n1684 ), .Y(\U1/aes_core/SB3/n3208 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1674  ( .A(\U1/aes_core/SB3/n3208 ), .Y(
        \U1/aes_core/SB3/n3194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1673  ( .A(\U1/aes_core/SB3/n1030 ), .B(
        Dout[4]), .Y(\U1/aes_core/SB3/n1708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1672  ( .A(\U1/aes_core/SB3/n1700 ), .B(
        \U1/aes_core/SB3/n1708 ), .Y(\U1/aes_core/SB3/n3248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1671  ( .A(\U1/aes_core/SB3/n3096 ), .B(
        \U1/aes_core/SB3/n3248 ), .Y(\U1/aes_core/SB3/n2987 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1670  ( .A(\U1/aes_core/SB3/n1203 ), .B(
        \U1/aes_core/SB3/n1158 ), .Y(\U1/aes_core/SB3/n1699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1669  ( .A(\U1/aes_core/SB3/n1690 ), .B(
        \U1/aes_core/SB3/n1699 ), .Y(\U1/aes_core/SB3/n3223 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1668  ( .A(\U1/aes_core/SB3/n3223 ), .Y(
        \U1/aes_core/SB3/n2968 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1667  ( .A0(\U1/aes_core/SB3/n3194 ), 
        .A1(\U1/aes_core/SB3/n2987 ), .B0(\U1/aes_core/SB3/n2968 ), .B1(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n1218 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1666  ( .AN(\U1/aes_core/SB3/n3009 ), 
        .B(\U1/aes_core/SB3/n1621 ), .C(\U1/aes_core/SB3/n1218 ), .Y(
        \U1/aes_core/SB3/n1721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1665  ( .A(\U1/aes_core/SB3/n1682 ), .B(
        \U1/aes_core/SB3/n1699 ), .Y(\U1/aes_core/SB3/n3113 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1664  ( .A(\U1/aes_core/SB3/n1686 ), .B(
        \U1/aes_core/SB3/n1687 ), .Y(\U1/aes_core/SB3/n3258 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1663  ( .A(\U1/aes_core/SB3/n1709 ), .B(
        \U1/aes_core/SB3/n1690 ), .Y(\U1/aes_core/SB3/n3164 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1662  ( .A(\U1/aes_core/SB3/n1686 ), .B(
        \U1/aes_core/SB3/n1692 ), .Y(\U1/aes_core/SB3/n3161 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1661  ( .A(\U1/aes_core/SB3/n1683 ), .B(
        \U1/aes_core/SB3/n1693 ), .Y(\U1/aes_core/SB3/n3166 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1660  ( .A(\U1/aes_core/SB3/n3166 ), .Y(
        \U1/aes_core/SB3/n3146 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1659  ( .A(\U1/aes_core/SB3/n3248 ), .Y(
        \U1/aes_core/SB3/n2982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1658  ( .A(\U1/aes_core/SB3/n1684 ), .B(
        \U1/aes_core/SB3/n1692 ), .Y(\U1/aes_core/SB3/n3184 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1657  ( .A(\U1/aes_core/SB3/n3184 ), .Y(
        \U1/aes_core/SB3/n3209 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1656  ( .A0(\U1/aes_core/SB3/n3146 ), 
        .A1(\U1/aes_core/SB3/n3210 ), .B0(\U1/aes_core/SB3/n2982 ), .B1(
        \U1/aes_core/SB3/n3209 ), .Y(\U1/aes_core/SB3/n1685 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1655  ( .A0(\U1/aes_core/SB3/n3113 ), 
        .A1(\U1/aes_core/SB3/n3258 ), .B0(\U1/aes_core/SB3/n3164 ), .B1(
        \U1/aes_core/SB3/n3161 ), .C0(\U1/aes_core/SB3/n1685 ), .Y(
        \U1/aes_core/SB3/n1720 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1654  ( .A(\U1/aes_core/SB3/n3166 ), .B(
        \U1/aes_core/SB3/n3113 ), .Y(\U1/aes_core/SB3/n2975 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1653  ( .A(\U1/aes_core/SB3/n3161 ), .B(
        \U1/aes_core/SB3/n3096 ), .Y(\U1/aes_core/SB3/n2985 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1652  ( .A(\U1/aes_core/SB3/n2985 ), .Y(
        \U1/aes_core/SB3/n1689 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1651  ( .A(\U1/aes_core/SB3/n1686 ), .B(
        \U1/aes_core/SB3/n1702 ), .Y(\U1/aes_core/SB3/n3236 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1650  ( .A(\U1/aes_core/SB3/n3236 ), .Y(
        \U1/aes_core/SB3/n3185 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1649  ( .A(\U1/aes_core/SB3/n1687 ), .B(
        \U1/aes_core/SB3/n1693 ), .Y(\U1/aes_core/SB3/n3221 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1648  ( .A(\U1/aes_core/SB3/n3221 ), .Y(
        \U1/aes_core/SB3/n3232 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1647  ( .A0(\U1/aes_core/SB3/n3185 ), 
        .A1(\U1/aes_core/SB3/n3232 ), .B0(\U1/aes_core/SB3/n3186 ), .Y(
        \U1/aes_core/SB3/n1688 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1646  ( .A(\U1/aes_core/SB3/n1691 ), .B(
        \U1/aes_core/SB3/n1708 ), .Y(\U1/aes_core/SB3/n3237 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1645  ( .A(\U1/aes_core/SB3/n3237 ), .Y(
        \U1/aes_core/SB3/n3187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1644  ( .A(\U1/aes_core/SB3/n3187 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3002 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1643  ( .AN(\U1/aes_core/SB3/n2975 ), 
        .B(\U1/aes_core/SB3/n1689 ), .C(\U1/aes_core/SB3/n1688 ), .D(
        \U1/aes_core/SB3/n3002 ), .Y(\U1/aes_core/SB3/n1698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1642  ( .A(\U1/aes_core/SB3/n1701 ), .B(
        \U1/aes_core/SB3/n1699 ), .Y(\U1/aes_core/SB3/n3257 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1641  ( .A(\U1/aes_core/SB3/n1691 ), .B(
        \U1/aes_core/SB3/n1690 ), .Y(\U1/aes_core/SB3/n3249 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1640  ( .A0(\U1/aes_core/SB3/n2327 ), 
        .A1(\U1/aes_core/SB3/n3076 ), .B0(\U1/aes_core/SB3/n3257 ), .B1(
        \U1/aes_core/SB3/n3166 ), .C0(\U1/aes_core/SB3/n3249 ), .C1(
        \U1/aes_core/SB3/n3184 ), .Y(\U1/aes_core/SB3/n1697 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1639  ( .A(\U1/aes_core/SB3/n3208 ), .B(
        \U1/aes_core/SB3/n2327 ), .Y(\U1/aes_core/SB3/n3060 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1638  ( .A(\U1/aes_core/SB3/n2982 ), .B(
        \U1/aes_core/SB3/n3146 ), .Y(\U1/aes_core/SB3/n3013 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1637  ( .A(\U1/aes_core/SB3/n3209 ), .B(
        \U1/aes_core/SB3/n3210 ), .Y(\U1/aes_core/SB3/n3033 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1636  ( .A(\U1/aes_core/SB3/n3164 ), .Y(
        \U1/aes_core/SB3/n3238 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1635  ( .A(\U1/aes_core/SB3/n3238 ), .B(
        \U1/aes_core/SB3/n3068 ), .Y(\U1/aes_core/SB3/n3071 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1634  ( .AN(\U1/aes_core/SB3/n3060 ), 
        .B(\U1/aes_core/SB3/n3013 ), .C(\U1/aes_core/SB3/n3033 ), .D(
        \U1/aes_core/SB3/n3071 ), .Y(\U1/aes_core/SB3/n1696 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1633  ( .A(\U1/aes_core/SB3/n1709 ), .B(
        \U1/aes_core/SB3/n1701 ), .Y(\U1/aes_core/SB3/n2983 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1632  ( .A(\U1/aes_core/SB3/n2983 ), .B(
        \U1/aes_core/SB3/n3220 ), .Y(\U1/aes_core/SB3/n3137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1631  ( .A(\U1/aes_core/SB3/n1693 ), .B(
        \U1/aes_core/SB3/n1692 ), .Y(\U1/aes_core/SB3/n3256 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1630  ( .A(\U1/aes_core/SB3/n3223 ), .B(
        \U1/aes_core/SB3/n3256 ), .Y(\U1/aes_core/SB3/n3102 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1629  ( .A(\U1/aes_core/SB3/n3102 ), .Y(
        \U1/aes_core/SB3/n1694 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1628  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3068 ), .Y(\U1/aes_core/SB3/n3121 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1627  ( .A(\U1/aes_core/SB3/n3256 ), .Y(
        \U1/aes_core/SB3/n3239 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1626  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3239 ), .Y(\U1/aes_core/SB3/n3172 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1625  ( .AN(\U1/aes_core/SB3/n3137 ), 
        .B(\U1/aes_core/SB3/n1694 ), .C(\U1/aes_core/SB3/n3121 ), .D(
        \U1/aes_core/SB3/n3172 ), .Y(\U1/aes_core/SB3/n1695 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1624  ( .A(\U1/aes_core/SB3/n1698 ), .B(
        \U1/aes_core/SB3/n1697 ), .C(\U1/aes_core/SB3/n1696 ), .D(
        \U1/aes_core/SB3/n1695 ), .Y(\U1/aes_core/SB3/n2905 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1623  ( .A(\U1/aes_core/SB3/n3163 ), .B(
        \U1/aes_core/SB3/n2983 ), .Y(\U1/aes_core/SB3/n3171 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1622  ( .A(\U1/aes_core/SB3/n1708 ), .B(
        \U1/aes_core/SB3/n1699 ), .Y(\U1/aes_core/SB3/n3079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1621  ( .A(\U1/aes_core/SB3/n3145 ), .B(
        \U1/aes_core/SB3/n3079 ), .Y(\U1/aes_core/SB3/n3050 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1620  ( .A(\U1/aes_core/SB3/n3257 ), .Y(
        \U1/aes_core/SB3/n3213 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1619  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3194 ), .Y(\U1/aes_core/SB3/n2999 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1618  ( .A0(\U1/aes_core/SB3/n3079 ), 
        .A1(\U1/aes_core/SB3/n3256 ), .B0(\U1/aes_core/SB3/n2999 ), .Y(
        \U1/aes_core/SB3/n1707 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1617  ( .A(\U1/aes_core/SB3/n3094 ), .Y(
        \U1/aes_core/SB3/n3189 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1616  ( .A(\U1/aes_core/SB3/n3189 ), .B(
        \U1/aes_core/SB3/n3212 ), .Y(\U1/aes_core/SB3/n3190 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1615  ( .A(\U1/aes_core/SB3/n3212 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1614  ( .A(\U1/aes_core/SB3/n1701 ), .B(
        \U1/aes_core/SB3/n1700 ), .Y(\U1/aes_core/SB3/n3219 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1613  ( .A(\U1/aes_core/SB3/n3219 ), .Y(
        \U1/aes_core/SB3/n2994 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1612  ( .A(\U1/aes_core/SB3/n3185 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3018 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1611  ( .A(\U1/aes_core/SB3/n3207 ), .Y(
        \U1/aes_core/SB3/n3188 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1610  ( .A(\U1/aes_core/SB3/n3188 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3082 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1609  ( .A(\U1/aes_core/SB3/n3190 ), .B(
        \U1/aes_core/SB3/n3149 ), .C(\U1/aes_core/SB3/n3018 ), .D(
        \U1/aes_core/SB3/n3082 ), .Y(\U1/aes_core/SB3/n1706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1608  ( .A(\U1/aes_core/SB3/n3209 ), .B(
        \U1/aes_core/SB3/n3187 ), .Y(\U1/aes_core/SB3/n3116 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1607  ( .A(\U1/aes_core/SB3/n3251 ), .B(
        \U1/aes_core/SB3/n3187 ), .Y(\U1/aes_core/SB3/n3107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1606  ( .A(\U1/aes_core/SB3/n3249 ), .Y(
        \U1/aes_core/SB3/n3242 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1605  ( .A(\U1/aes_core/SB3/n3146 ), .B(
        \U1/aes_core/SB3/n3242 ), .Y(\U1/aes_core/SB3/n2979 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1604  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3185 ), .Y(\U1/aes_core/SB3/n3090 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1603  ( .A(\U1/aes_core/SB3/n3116 ), .B(
        \U1/aes_core/SB3/n3107 ), .C(\U1/aes_core/SB3/n2979 ), .D(
        \U1/aes_core/SB3/n3090 ), .Y(\U1/aes_core/SB3/n1705 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1602  ( .A(\U1/aes_core/SB3/n3161 ), .Y(
        \U1/aes_core/SB3/n3130 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1601  ( .A(\U1/aes_core/SB3/n2982 ), .B(
        \U1/aes_core/SB3/n3130 ), .Y(\U1/aes_core/SB3/n2966 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1600  ( .A(\U1/aes_core/SB3/n1703 ), .B(
        \U1/aes_core/SB3/n1702 ), .Y(\U1/aes_core/SB3/n3196 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1599  ( .A(\U1/aes_core/SB3/n3196 ), .Y(
        \U1/aes_core/SB3/n3230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1598  ( .A(\U1/aes_core/SB3/n2982 ), .B(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n3030 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1597  ( .A(\U1/aes_core/SB3/n3145 ), .Y(
        \U1/aes_core/SB3/n3253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1596  ( .A(\U1/aes_core/SB3/n3253 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n3065 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1595  ( .A(\U1/aes_core/SB3/n3186 ), .B(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n3214 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1594  ( .A(\U1/aes_core/SB3/n2966 ), .B(
        \U1/aes_core/SB3/n3030 ), .C(\U1/aes_core/SB3/n3065 ), .D(
        \U1/aes_core/SB3/n3214 ), .Y(\U1/aes_core/SB3/n1704 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1593  ( .A(\U1/aes_core/SB3/n3171 ), .B(
        \U1/aes_core/SB3/n3050 ), .C(\U1/aes_core/SB3/n1707 ), .D(
        \U1/aes_core/SB3/n1706 ), .E(\U1/aes_core/SB3/n1705 ), .F(
        \U1/aes_core/SB3/n1704 ), .Y(\U1/aes_core/SB3/n2894 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1592  ( .A(\U1/aes_core/SB3/n2894 ), .Y(
        \U1/aes_core/SB3/n1718 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1591  ( .A(\U1/aes_core/SB3/n3221 ), .B(
        \U1/aes_core/SB3/n3079 ), .Y(\U1/aes_core/SB3/n2976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1590  ( .A(\U1/aes_core/SB3/n1709 ), .B(
        \U1/aes_core/SB3/n1708 ), .Y(\U1/aes_core/SB3/n3218 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1589  ( .A(\U1/aes_core/SB3/n3218 ), .B(
        \U1/aes_core/SB3/n3094 ), .Y(\U1/aes_core/SB3/n3103 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1588  ( .A(\U1/aes_core/SB3/n3103 ), .Y(
        \U1/aes_core/SB3/n1711 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1587  ( .A(\U1/aes_core/SB3/n3096 ), .Y(
        \U1/aes_core/SB3/n3243 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1586  ( .A0(\U1/aes_core/SB3/n2994 ), 
        .A1(\U1/aes_core/SB3/n3243 ), .B0(\U1/aes_core/SB3/n3230 ), .Y(
        \U1/aes_core/SB3/n1710 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1585  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3130 ), .Y(\U1/aes_core/SB3/n3001 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1584  ( .AN(\U1/aes_core/SB3/n2976 ), 
        .B(\U1/aes_core/SB3/n1711 ), .C(\U1/aes_core/SB3/n1710 ), .D(
        \U1/aes_core/SB3/n3001 ), .Y(\U1/aes_core/SB3/n1715 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1583  ( .A0(\U1/aes_core/SB3/n3207 ), 
        .A1(\U1/aes_core/SB3/n3255 ), .B0(\U1/aes_core/SB3/n3113 ), .B1(
        \U1/aes_core/SB3/n3161 ), .C0(\U1/aes_core/SB3/n3220 ), .C1(
        \U1/aes_core/SB3/n3237 ), .Y(\U1/aes_core/SB3/n1714 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1582  ( .A(\U1/aes_core/SB3/n3255 ), .B(
        \U1/aes_core/SB3/n3258 ), .Y(\U1/aes_core/SB3/n3041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1581  ( .A(\U1/aes_core/SB3/n3243 ), .B(
        \U1/aes_core/SB3/n3185 ), .Y(\U1/aes_core/SB3/n3174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1580  ( .A(\U1/aes_core/SB3/n3146 ), .B(
        \U1/aes_core/SB3/n3243 ), .Y(\U1/aes_core/SB3/n3108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1579  ( .A(\U1/aes_core/SB3/n3130 ), .B(
        \U1/aes_core/SB3/n3210 ), .Y(\U1/aes_core/SB3/n2980 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1578  ( .AN(\U1/aes_core/SB3/n3041 ), 
        .B(\U1/aes_core/SB3/n3174 ), .C(\U1/aes_core/SB3/n3108 ), .D(
        \U1/aes_core/SB3/n2980 ), .Y(\U1/aes_core/SB3/n1713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1577  ( .A(\U1/aes_core/SB3/n3253 ), .B(
        \U1/aes_core/SB3/n3238 ), .Y(\U1/aes_core/SB3/n3053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1576  ( .A(\U1/aes_core/SB3/n3130 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3120 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1575  ( .A(\U1/aes_core/SB3/n2982 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3021 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1574  ( .A(\U1/aes_core/SB3/n3189 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n3066 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1573  ( .A(\U1/aes_core/SB3/n3053 ), .B(
        \U1/aes_core/SB3/n3120 ), .C(\U1/aes_core/SB3/n3021 ), .D(
        \U1/aes_core/SB3/n3066 ), .Y(\U1/aes_core/SB3/n1712 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1572  ( .A(\U1/aes_core/SB3/n1715 ), .B(
        \U1/aes_core/SB3/n1714 ), .C(\U1/aes_core/SB3/n1713 ), .D(
        \U1/aes_core/SB3/n1712 ), .Y(\U1/aes_core/SB3/n1716 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1571  ( .A(\U1/aes_core/SB3/n1716 ), .Y(
        \U1/aes_core/SB3/n3235 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1570  ( .A(\U1/aes_core/SB3/n3251 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n1717 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1569  ( .AN(\U1/aes_core/SB3/n2905 ), 
        .B(\U1/aes_core/SB3/n1718 ), .C(\U1/aes_core/SB3/n3235 ), .D(
        \U1/aes_core/SB3/n1717 ), .Y(\U1/aes_core/SB3/n1719 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1568  ( .A(\U1/aes_core/SB3/n3014 ), .B(
        \U1/aes_core/SB3/n3111 ), .C(\U1/aes_core/SB3/n1722 ), .D(
        \U1/aes_core/SB3/n1721 ), .E(\U1/aes_core/SB3/n1720 ), .F(
        \U1/aes_core/SB3/n1719 ), .Y(\U1/aes_core/SB3/n2346 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1567  ( .A(\U1/aes_core/SB3/n3236 ), .B(
        \U1/aes_core/SB3/n2327 ), .Y(\U1/aes_core/SB3/n3059 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1566  ( .A(\U1/aes_core/SB3/n3186 ), .B(
        \U1/aes_core/SB3/n3253 ), .Y(\U1/aes_core/SB3/n3110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1565  ( .A(\U1/aes_core/SB3/n3242 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3012 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1564  ( .A(\U1/aes_core/SB3/n2983 ), .Y(
        \U1/aes_core/SB3/n3231 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1563  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3035 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1562  ( .AN(\U1/aes_core/SB3/n3059 ), 
        .B(\U1/aes_core/SB3/n3110 ), .C(\U1/aes_core/SB3/n3012 ), .D(
        \U1/aes_core/SB3/n3035 ), .Y(\U1/aes_core/SB3/n1729 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1561  ( .A(\U1/aes_core/SB3/n3223 ), .B(
        \U1/aes_core/SB3/n3094 ), .Y(\U1/aes_core/SB3/n3136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1560  ( .A(\U1/aes_core/SB3/n3146 ), .B(
        \U1/aes_core/SB3/n3212 ), .Y(\U1/aes_core/SB3/n2992 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1559  ( .A0(\U1/aes_core/SB3/n3232 ), 
        .A1(\U1/aes_core/SB3/n3152 ), .B0(\U1/aes_core/SB3/n2982 ), .Y(
        \U1/aes_core/SB3/n1723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1558  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3084 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1557  ( .AN(\U1/aes_core/SB3/n3136 ), 
        .B(\U1/aes_core/SB3/n2992 ), .C(\U1/aes_core/SB3/n1723 ), .D(
        \U1/aes_core/SB3/n3084 ), .Y(\U1/aes_core/SB3/n1724 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1556  ( .A(\U1/aes_core/SB3/n1724 ), .Y(
        \U1/aes_core/SB3/n1728 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1555  ( .A(\U1/aes_core/SB3/n3113 ), .Y(
        \U1/aes_core/SB3/n3233 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1554  ( .A(\U1/aes_core/SB3/n3258 ), .Y(
        \U1/aes_core/SB3/n3153 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U1553  ( .A0(\U1/aes_core/SB3/n3253 ), 
        .A1(\U1/aes_core/SB3/n3187 ), .B0(\U1/aes_core/SB3/n3233 ), .B1(
        \U1/aes_core/SB3/n3068 ), .C0(\U1/aes_core/SB3/n3153 ), .C1(
        \U1/aes_core/SB3/n3231 ), .Y(\U1/aes_core/SB3/n1727 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1552  ( .A0(\U1/aes_core/SB3/n3079 ), 
        .A1(\U1/aes_core/SB3/n3236 ), .B0(\U1/aes_core/SB3/n3256 ), .B1(
        \U1/aes_core/SB3/n3257 ), .Y(\U1/aes_core/SB3/n1725 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1551  ( .A0(\U1/aes_core/SB3/n3130 ), 
        .A1(\U1/aes_core/SB3/n2968 ), .B0(\U1/aes_core/SB3/n3186 ), .B1(
        \U1/aes_core/SB3/n3209 ), .C0(\U1/aes_core/SB3/n1725 ), .Y(
        \U1/aes_core/SB3/n1726 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1550  ( .AN(\U1/aes_core/SB3/n1729 ), 
        .B(\U1/aes_core/SB3/n1728 ), .C(\U1/aes_core/SB3/n1727 ), .D(
        \U1/aes_core/SB3/n1726 ), .Y(\U1/aes_core/SB3/n2903 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1549  ( .A(\U1/aes_core/SB3/n3257 ), .B(
        \U1/aes_core/SB3/n3094 ), .Y(\U1/aes_core/SB3/n2977 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1548  ( .A0(\U1/aes_core/SB3/n3164 ), 
        .A1(\U1/aes_core/SB3/n3257 ), .B0(\U1/aes_core/SB3/n3196 ), .Y(
        \U1/aes_core/SB3/n1734 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1547  ( .A(\U1/aes_core/SB3/n3196 ), .B(
        \U1/aes_core/SB3/n3184 ), .Y(\U1/aes_core/SB3/n3061 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB3/U1546  ( .A0(\U1/aes_core/SB3/n3185 ), 
        .A1(\U1/aes_core/SB3/n2968 ), .B0(\U1/aes_core/SB3/n3061 ), .B1(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n1733 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1545  ( .A0(\U1/aes_core/SB3/n3218 ), 
        .A1(\U1/aes_core/SB3/n3258 ), .B0(\U1/aes_core/SB3/n2983 ), .B1(
        \U1/aes_core/SB3/n3076 ), .C0(\U1/aes_core/SB3/n3220 ), .C1(
        \U1/aes_core/SB3/n3249 ), .Y(\U1/aes_core/SB3/n1732 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1544  ( .A(\U1/aes_core/SB3/n3079 ), .Y(
        \U1/aes_core/SB3/n3147 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1543  ( .A(\U1/aes_core/SB3/n3251 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3173 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1542  ( .A(\U1/aes_core/SB3/n3146 ), .B(
        \U1/aes_core/SB3/n2968 ), .Y(\U1/aes_core/SB3/n3000 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1541  ( .A(\U1/aes_core/SB3/n2982 ), .B(
        \U1/aes_core/SB3/n3189 ), .Y(\U1/aes_core/SB3/n3020 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1540  ( .A(\U1/aes_core/SB3/n3146 ), .B(
        \U1/aes_core/SB3/n3187 ), .Y(\U1/aes_core/SB3/n3119 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1539  ( .A(\U1/aes_core/SB3/n3173 ), .B(
        \U1/aes_core/SB3/n3000 ), .C(\U1/aes_core/SB3/n3020 ), .D(
        \U1/aes_core/SB3/n3119 ), .Y(\U1/aes_core/SB3/n1731 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1538  ( .A(\U1/aes_core/SB3/n3166 ), .B(
        \U1/aes_core/SB3/n3079 ), .Y(\U1/aes_core/SB3/n3042 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1537  ( .A(\U1/aes_core/SB3/n3152 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3052 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1536  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3068 ), .Y(\U1/aes_core/SB3/n3083 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1535  ( .AN(\U1/aes_core/SB3/n3042 ), 
        .B(\U1/aes_core/SB3/n3052 ), .C(\U1/aes_core/SB3/n3083 ), .Y(
        \U1/aes_core/SB3/n1730 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1534  ( .A(\U1/aes_core/SB3/n2977 ), .B(
        \U1/aes_core/SB3/n1734 ), .C(\U1/aes_core/SB3/n1733 ), .D(
        \U1/aes_core/SB3/n1732 ), .E(\U1/aes_core/SB3/n1731 ), .F(
        \U1/aes_core/SB3/n1730 ), .Y(\U1/aes_core/SB3/n3264 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1533  ( .A0(\U1/aes_core/SB3/n2982 ), 
        .A1(\U1/aes_core/SB3/n3210 ), .B0(\U1/aes_core/SB3/n3241 ), .Y(
        \U1/aes_core/SB3/n1735 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1532  ( .A(\U1/aes_core/SB3/n2968 ), .B(
        \U1/aes_core/SB3/n3068 ), .Y(\U1/aes_core/SB3/n3105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1531  ( .A(\U1/aes_core/SB3/n3185 ), .B(
        \U1/aes_core/SB3/n3233 ), .Y(\U1/aes_core/SB3/n2997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1530  ( .A(\U1/aes_core/SB3/n3233 ), .B(
        \U1/aes_core/SB3/n3189 ), .Y(\U1/aes_core/SB3/n3048 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1529  ( .A(\U1/aes_core/SB3/n1735 ), .B(
        \U1/aes_core/SB3/n3105 ), .C(\U1/aes_core/SB3/n2997 ), .D(
        \U1/aes_core/SB3/n3048 ), .Y(\U1/aes_core/SB3/n1739 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1528  ( .A0(\U1/aes_core/SB3/n3236 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n2983 ), .B1(
        \U1/aes_core/SB3/n3208 ), .C0(\U1/aes_core/SB3/n3237 ), .C1(
        \U1/aes_core/SB3/n3094 ), .Y(\U1/aes_core/SB3/n1738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1527  ( .A(\U1/aes_core/SB3/n3188 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n3029 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1526  ( .A(\U1/aes_core/SB3/n3187 ), .B(
        \U1/aes_core/SB3/n3239 ), .Y(\U1/aes_core/SB3/n3169 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1525  ( .A(\U1/aes_core/SB3/n3187 ), .B(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n3016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1524  ( .A(\U1/aes_core/SB3/n3242 ), .B(
        \U1/aes_core/SB3/n3232 ), .Y(\U1/aes_core/SB3/n2978 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1523  ( .A(\U1/aes_core/SB3/n3029 ), .B(
        \U1/aes_core/SB3/n3169 ), .C(\U1/aes_core/SB3/n3016 ), .D(
        \U1/aes_core/SB3/n2978 ), .Y(\U1/aes_core/SB3/n1737 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1522  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1521  ( .A(\U1/aes_core/SB3/n3251 ), .B(
        \U1/aes_core/SB3/n3212 ), .Y(\U1/aes_core/SB3/n3064 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1520  ( .A(\U1/aes_core/SB3/n3241 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1519  ( .A(\U1/aes_core/SB3/n2994 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n2965 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1518  ( .A(\U1/aes_core/SB3/n3091 ), .B(
        \U1/aes_core/SB3/n3064 ), .C(\U1/aes_core/SB3/n3115 ), .D(
        \U1/aes_core/SB3/n2965 ), .Y(\U1/aes_core/SB3/n1736 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1517  ( .A(\U1/aes_core/SB3/n1739 ), .B(
        \U1/aes_core/SB3/n1738 ), .C(\U1/aes_core/SB3/n1737 ), .D(
        \U1/aes_core/SB3/n1736 ), .Y(\U1/aes_core/SB3/n2892 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1516  ( .A(\U1/aes_core/SB3/n2346 ), .B(
        \U1/aes_core/SB3/n2903 ), .C(\U1/aes_core/SB3/n3264 ), .D(
        \U1/aes_core/SB3/n2892 ), .Y(\U1/aes_core/SB3/n1748 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1515  ( .A(\U1/aes_core/SB3/n3218 ), .Y(
        \U1/aes_core/SB3/n3142 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1514  ( .A0(\U1/aes_core/SB3/n3094 ), 
        .A1(\U1/aes_core/SB3/n2328 ), .B0(\U1/aes_core/SB3/n3063 ), .B1(
        \U1/aes_core/SB3/n3249 ), .Y(\U1/aes_core/SB3/n1740 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1513  ( .A0(\U1/aes_core/SB3/n3142 ), 
        .A1(\U1/aes_core/SB3/n3194 ), .B0(\U1/aes_core/SB3/n3243 ), .B1(
        \U1/aes_core/SB3/n3251 ), .C0(\U1/aes_core/SB3/n1740 ), .Y(
        \U1/aes_core/SB3/n1747 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1512  ( .A(\U1/aes_core/SB3/n3163 ), .B(
        \U1/aes_core/SB3/n3166 ), .Y(\U1/aes_core/SB3/n3162 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1511  ( .A0(\U1/aes_core/SB3/n3097 ), 
        .A1(\U1/aes_core/SB3/n3166 ), .B0(\U1/aes_core/SB3/n3079 ), .B1(
        \U1/aes_core/SB3/n3207 ), .Y(\U1/aes_core/SB3/n1741 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1510  ( .A0(\U1/aes_core/SB3/n2994 ), 
        .A1(\U1/aes_core/SB3/n3162 ), .B0(\U1/aes_core/SB3/n3213 ), .B1(
        \U1/aes_core/SB3/n3232 ), .C0(\U1/aes_core/SB3/n1741 ), .Y(
        \U1/aes_core/SB3/n1746 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1509  ( .A(\U1/aes_core/SB3/n3237 ), .B(
        \U1/aes_core/SB3/n3096 ), .Y(\U1/aes_core/SB3/n1744 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1508  ( .A(\U1/aes_core/SB3/n3187 ), .B(
        \U1/aes_core/SB3/n3212 ), .Y(\U1/aes_core/SB3/n3154 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1507  ( .A(\U1/aes_core/SB3/n3154 ), .Y(
        \U1/aes_core/SB3/n1743 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1506  ( .A(\U1/aes_core/SB3/n3145 ), .B(
        \U1/aes_core/SB3/n3218 ), .Y(\U1/aes_core/SB3/n3026 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1505  ( .A(\U1/aes_core/SB3/n3223 ), .B(
        \U1/aes_core/SB3/n3221 ), .Y(\U1/aes_core/SB3/n3179 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1503  ( .A(\U1/aes_core/SB3/n3194 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3036 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1501  ( .A0(\U1/aes_core/SB3/n3153 ), 
        .A1(\U1/aes_core/SB3/n1744 ), .B0(\U1/aes_core/SB3/n3130 ), .B1(
        \U1/aes_core/SB3/n1743 ), .C0(\U1/aes_core/SB3/n1742 ), .Y(
        \U1/aes_core/SB3/n1745 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1500  ( .AN(\U1/aes_core/SB3/n1748 ), 
        .B(\U1/aes_core/SB3/n1747 ), .C(\U1/aes_core/SB3/n1746 ), .D(
        \U1/aes_core/SB3/n1745 ), .Y(\U1/aes_core/sb3 [0]) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1499  ( .A(Dout[14]), .Y(
        \U1/aes_core/SB3/n1755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1498  ( .A(Dout[15]), .Y(
        \U1/aes_core/SB3/n1750 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1497  ( .A(\U1/aes_core/SB3/n1755 ), .B(
        \U1/aes_core/SB3/n1750 ), .Y(\U1/aes_core/SB3/n1760 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1496  ( .A(Dout[13]), .Y(
        \U1/aes_core/SB3/n1749 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1495  ( .A(\U1/aes_core/SB3/n1749 ), .B(
        Dout[12]), .Y(\U1/aes_core/SB3/n1767 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1494  ( .A(\U1/aes_core/SB3/n1760 ), .B(
        \U1/aes_core/SB3/n1767 ), .Y(\U1/aes_core/SB3/n3300 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1493  ( .A(Dout[11]), .Y(
        \U1/aes_core/SB3/n1758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1492  ( .A(\U1/aes_core/SB3/n1758 ), .B(
        Dout[10]), .Y(\U1/aes_core/SB3/n1773 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1491  ( .A(Dout[8]), .Y(
        \U1/aes_core/SB3/n1751 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1490  ( .A(\U1/aes_core/SB3/n1751 ), .B(
        Dout[9]), .Y(\U1/aes_core/SB3/n1761 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1489  ( .A(\U1/aes_core/SB3/n1773 ), .B(
        \U1/aes_core/SB3/n1761 ), .Y(\U1/aes_core/SB3/n1912 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1488  ( .A(\U1/aes_core/SB3/n3300 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n1821 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1487  ( .A(Dout[9]), .Y(
        \U1/aes_core/SB3/n1752 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1486  ( .A(\U1/aes_core/SB3/n1752 ), .B(
        Dout[8]), .Y(\U1/aes_core/SB3/n1770 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1485  ( .A(Dout[10]), .Y(
        \U1/aes_core/SB3/n1757 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1484  ( .A(\U1/aes_core/SB3/n1757 ), .B(
        Dout[11]), .Y(\U1/aes_core/SB3/n1754 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1483  ( .A(\U1/aes_core/SB3/n1770 ), .B(
        \U1/aes_core/SB3/n1754 ), .Y(\U1/aes_core/SB3/n3346 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1482  ( .A(Dout[12]), .Y(
        \U1/aes_core/SB3/n1753 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1481  ( .A(\U1/aes_core/SB3/n1749 ), .B(
        \U1/aes_core/SB3/n1753 ), .Y(\U1/aes_core/SB3/n1781 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1480  ( .A(\U1/aes_core/SB3/n1750 ), .B(
        Dout[14]), .Y(\U1/aes_core/SB3/n1756 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1479  ( .A(\U1/aes_core/SB3/n1781 ), .B(
        \U1/aes_core/SB3/n1756 ), .Y(\U1/aes_core/SB3/n2021 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1478  ( .A0(\U1/aes_core/SB3/n1912 ), 
        .A1(\U1/aes_core/SB3/n3346 ), .B0(\U1/aes_core/SB3/n2021 ), .Y(
        \U1/aes_core/SB3/n1766 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1477  ( .A(\U1/aes_core/SB3/n1752 ), .B(
        \U1/aes_core/SB3/n1751 ), .Y(\U1/aes_core/SB3/n1772 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1476  ( .A(\U1/aes_core/SB3/n1754 ), .B(
        \U1/aes_core/SB3/n1772 ), .Y(\U1/aes_core/SB3/n2020 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1475  ( .A(\U1/aes_core/SB3/n1753 ), .B(
        Dout[13]), .Y(\U1/aes_core/SB3/n1783 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1474  ( .A(\U1/aes_core/SB3/n1760 ), .B(
        \U1/aes_core/SB3/n1783 ), .Y(\U1/aes_core/SB3/n1995 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1473  ( .A(Dout[11]), .B(Dout[10]), .Y(
        \U1/aes_core/SB3/n1780 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1472  ( .A(\U1/aes_core/SB3/n1772 ), .B(
        \U1/aes_core/SB3/n1780 ), .Y(\U1/aes_core/SB3/n3301 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1471  ( .A(\U1/aes_core/SB3/n3301 ), .Y(
        \U1/aes_core/SB3/n3339 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1470  ( .A(Dout[9]), .B(Dout[8]), .Y(
        \U1/aes_core/SB3/n1779 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1469  ( .A(\U1/aes_core/SB3/n1754 ), .B(
        \U1/aes_core/SB3/n1779 ), .Y(\U1/aes_core/SB3/n3296 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1468  ( .A(\U1/aes_core/SB3/n3296 ), .Y(
        \U1/aes_core/SB3/n3333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1467  ( .A(\U1/aes_core/SB3/n3339 ), .B(
        \U1/aes_core/SB3/n3333 ), .Y(\U1/aes_core/SB3/n1823 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1466  ( .A(Dout[15]), .B(Dout[14]), .Y(
        \U1/aes_core/SB3/n1774 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1465  ( .A(\U1/aes_core/SB3/n1767 ), .B(
        \U1/aes_core/SB3/n1774 ), .Y(\U1/aes_core/SB3/n3309 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1464  ( .A0(\U1/aes_core/SB3/n2020 ), 
        .A1(\U1/aes_core/SB3/n1995 ), .B0(\U1/aes_core/SB3/n1823 ), .B1(
        \U1/aes_core/SB3/n3309 ), .Y(\U1/aes_core/SB3/n1765 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1463  ( .A(\U1/aes_core/SB3/n1754 ), .B(
        \U1/aes_core/SB3/n1761 ), .Y(\U1/aes_core/SB3/n1888 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1462  ( .A(\U1/aes_core/SB3/n1767 ), .B(
        \U1/aes_core/SB3/n1756 ), .Y(\U1/aes_core/SB3/n3344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1461  ( .A(Dout[13]), .B(Dout[12]), .Y(
        \U1/aes_core/SB3/n1759 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1460  ( .A(\U1/aes_core/SB3/n1760 ), .B(
        \U1/aes_core/SB3/n1759 ), .Y(\U1/aes_core/SB3/n3280 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1459  ( .A(\U1/aes_core/SB3/n1783 ), .B(
        \U1/aes_core/SB3/n1756 ), .Y(\U1/aes_core/SB3/n3278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1458  ( .A(\U1/aes_core/SB3/n1773 ), .B(
        \U1/aes_core/SB3/n1779 ), .Y(\U1/aes_core/SB3/n2010 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1457  ( .A0(\U1/aes_core/SB3/n1888 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n3301 ), .B1(
        \U1/aes_core/SB3/n3280 ), .C0(\U1/aes_core/SB3/n3278 ), .C1(
        \U1/aes_core/SB3/n2010 ), .Y(\U1/aes_core/SB3/n1764 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1456  ( .A(\U1/aes_core/SB3/n1755 ), .B(
        Dout[15]), .Y(\U1/aes_core/SB3/n1782 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1455  ( .A(\U1/aes_core/SB3/n1782 ), .B(
        \U1/aes_core/SB3/n1759 ), .Y(\U1/aes_core/SB3/n3308 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1454  ( .A(\U1/aes_core/SB3/n3308 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n1873 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1453  ( .A(\U1/aes_core/SB3/n1770 ), .B(
        \U1/aes_core/SB3/n1773 ), .Y(\U1/aes_core/SB3/n3342 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1452  ( .A(\U1/aes_core/SB3/n3342 ), .Y(
        \U1/aes_core/SB3/n2058 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1451  ( .A(\U1/aes_core/SB3/n1759 ), .B(
        \U1/aes_core/SB3/n1756 ), .Y(\U1/aes_core/SB3/n1806 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1450  ( .A(\U1/aes_core/SB3/n1806 ), .Y(
        \U1/aes_core/SB3/n3268 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1449  ( .A(\U1/aes_core/SB3/n2058 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n1856 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1448  ( .A(\U1/aes_core/SB3/n1758 ), .B(
        \U1/aes_core/SB3/n1757 ), .Y(\U1/aes_core/SB3/n1769 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1447  ( .A(\U1/aes_core/SB3/n1772 ), .B(
        \U1/aes_core/SB3/n1769 ), .Y(\U1/aes_core/SB3/n2006 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1446  ( .A(\U1/aes_core/SB3/n2006 ), .Y(
        \U1/aes_core/SB3/n2068 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U1445  ( .A(\U1/aes_core/SB3/n1774 ), .B(
        \U1/aes_core/SB3/n1759 ), .Y(\U1/aes_core/SB3/n3299 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1444  ( .A(\U1/aes_core/SB3/n2068 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1928 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1443  ( .A(\U1/aes_core/SB3/n1760 ), .B(
        \U1/aes_core/SB3/n1781 ), .Y(\U1/aes_core/SB3/n3347 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1442  ( .A(\U1/aes_core/SB3/n3347 ), .Y(
        \U1/aes_core/SB3/n3305 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1441  ( .A(\U1/aes_core/SB3/n3305 ), .B(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n1953 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1440  ( .AN(\U1/aes_core/SB3/n1873 ), 
        .B(\U1/aes_core/SB3/n1856 ), .C(\U1/aes_core/SB3/n1928 ), .D(
        \U1/aes_core/SB3/n1953 ), .Y(\U1/aes_core/SB3/n1763 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1439  ( .A(\U1/aes_core/SB3/n1995 ), .Y(
        \U1/aes_core/SB3/n3269 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1438  ( .A(\U1/aes_core/SB3/n1780 ), .B(
        \U1/aes_core/SB3/n1761 ), .Y(\U1/aes_core/SB3/n2017 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1437  ( .A(\U1/aes_core/SB3/n2017 ), .Y(
        \U1/aes_core/SB3/n2054 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1436  ( .A(\U1/aes_core/SB3/n3269 ), .B(
        \U1/aes_core/SB3/n2054 ), .Y(\U1/aes_core/SB3/n1843 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1435  ( .A(\U1/aes_core/SB3/n3278 ), .Y(
        \U1/aes_core/SB3/n3332 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1434  ( .A(\U1/aes_core/SB3/n1761 ), .B(
        \U1/aes_core/SB3/n1769 ), .Y(\U1/aes_core/SB3/n2057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1433  ( .A(\U1/aes_core/SB3/n2057 ), .Y(
        \U1/aes_core/SB3/n2019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1432  ( .A(\U1/aes_core/SB3/n3332 ), .B(
        \U1/aes_core/SB3/n2019 ), .Y(\U1/aes_core/SB3/n1879 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1431  ( .A(\U1/aes_core/SB3/n3269 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1966 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U1430  ( .A(\U1/aes_core/SB3/n1843 ), .B(
        \U1/aes_core/SB3/n1879 ), .C(\U1/aes_core/SB3/n1966 ), .Y(
        \U1/aes_core/SB3/n1762 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1429  ( .A(\U1/aes_core/SB3/n1821 ), .B(
        \U1/aes_core/SB3/n1766 ), .C(\U1/aes_core/SB3/n1765 ), .D(
        \U1/aes_core/SB3/n1764 ), .E(\U1/aes_core/SB3/n1763 ), .F(
        \U1/aes_core/SB3/n1762 ), .Y(\U1/aes_core/SB3/n3353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1428  ( .A(\U1/aes_core/SB3/n1995 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n1944 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1427  ( .A(\U1/aes_core/SB3/n2010 ), .Y(
        \U1/aes_core/SB3/n3330 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1426  ( .A(\U1/aes_core/SB3/n1888 ), .Y(
        \U1/aes_core/SB3/n3334 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1425  ( .A(\U1/aes_core/SB3/n1767 ), .B(
        \U1/aes_core/SB3/n1782 ), .Y(\U1/aes_core/SB3/n3343 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1424  ( .A(\U1/aes_core/SB3/n3343 ), .Y(
        \U1/aes_core/SB3/n3274 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1423  ( .A0(\U1/aes_core/SB3/n3330 ), 
        .A1(\U1/aes_core/SB3/n3334 ), .B0(\U1/aes_core/SB3/n3274 ), .Y(
        \U1/aes_core/SB3/n1768 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1422  ( .A(\U1/aes_core/SB3/n3305 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1903 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1421  ( .A(\U1/aes_core/SB3/n2021 ), .Y(
        \U1/aes_core/SB3/n2053 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1420  ( .A(\U1/aes_core/SB3/n3339 ), .B(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n1865 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1419  ( .AN(\U1/aes_core/SB3/n1944 ), 
        .B(\U1/aes_core/SB3/n1768 ), .C(\U1/aes_core/SB3/n1903 ), .D(
        \U1/aes_core/SB3/n1865 ), .Y(\U1/aes_core/SB3/n1778 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1418  ( .A(\U1/aes_core/SB3/n3309 ), .Y(
        \U1/aes_core/SB3/n1976 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1417  ( .A(\U1/aes_core/SB3/n1770 ), .B(
        \U1/aes_core/SB3/n1780 ), .Y(\U1/aes_core/SB3/n2039 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1416  ( .A(\U1/aes_core/SB3/n2039 ), .Y(
        \U1/aes_core/SB3/n3340 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1415  ( .A(\U1/aes_core/SB3/n3280 ), .Y(
        \U1/aes_core/SB3/n2055 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1414  ( .A(\U1/aes_core/SB3/n1779 ), .B(
        \U1/aes_core/SB3/n1769 ), .Y(\U1/aes_core/SB3/n3281 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1413  ( .A(\U1/aes_core/SB3/n3281 ), .Y(
        \U1/aes_core/SB3/n3331 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U1412  ( .A0(\U1/aes_core/SB3/n1976 ), 
        .A1(\U1/aes_core/SB3/n2068 ), .B0(\U1/aes_core/SB3/n3340 ), .B1(
        \U1/aes_core/SB3/n2055 ), .C0(\U1/aes_core/SB3/n3331 ), .C1(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n1777 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1411  ( .A(\U1/aes_core/SB3/n3300 ), .Y(
        \U1/aes_core/SB3/n1952 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1410  ( .A(\U1/aes_core/SB3/n1774 ), .B(
        \U1/aes_core/SB3/n1781 ), .Y(\U1/aes_core/SB3/n2070 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1409  ( .A(\U1/aes_core/SB3/n1770 ), .B(
        \U1/aes_core/SB3/n1769 ), .Y(\U1/aes_core/SB3/n3279 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1408  ( .A0(\U1/aes_core/SB3/n2070 ), 
        .A1(\U1/aes_core/SB3/n3346 ), .B0(\U1/aes_core/SB3/n3279 ), .B1(
        \U1/aes_core/SB3/n1995 ), .Y(\U1/aes_core/SB3/n1771 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1407  ( .A0(\U1/aes_core/SB3/n2058 ), 
        .A1(\U1/aes_core/SB3/n3305 ), .B0(\U1/aes_core/SB3/n1952 ), .B1(
        \U1/aes_core/SB3/n2019 ), .C0(\U1/aes_core/SB3/n1771 ), .Y(
        \U1/aes_core/SB3/n1776 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1406  ( .A(\U1/aes_core/SB3/n3268 ), .B(
        \U1/aes_core/SB3/n2019 ), .Y(\U1/aes_core/SB3/n1880 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1405  ( .A(\U1/aes_core/SB3/n1773 ), .B(
        \U1/aes_core/SB3/n1772 ), .Y(\U1/aes_core/SB3/n3302 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1404  ( .A(\U1/aes_core/SB3/n3302 ), .Y(
        \U1/aes_core/SB3/n3276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1403  ( .A(\U1/aes_core/SB3/n3276 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n1845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1402  ( .A(\U1/aes_core/SB3/n2070 ), .Y(
        \U1/aes_core/SB3/n3324 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1401  ( .A(\U1/aes_core/SB3/n3324 ), .B(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n1929 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1400  ( .A(\U1/aes_core/SB3/n1783 ), .B(
        \U1/aes_core/SB3/n1774 ), .Y(\U1/aes_core/SB3/n2065 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1399  ( .A(\U1/aes_core/SB3/n2065 ), .Y(
        \U1/aes_core/SB3/n3322 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1398  ( .A(\U1/aes_core/SB3/n3322 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1852 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB3/U1397  ( .A(\U1/aes_core/SB3/n1880 ), .B(
        \U1/aes_core/SB3/n1845 ), .C(\U1/aes_core/SB3/n1929 ), .D(
        \U1/aes_core/SB3/n1852 ), .Y(\U1/aes_core/SB3/n1775 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1396  ( .AN(\U1/aes_core/SB3/n1778 ), 
        .B(\U1/aes_core/SB3/n1777 ), .C(\U1/aes_core/SB3/n1776 ), .D(
        \U1/aes_core/SB3/n1775 ), .Y(\U1/aes_core/SB3/n3295 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1395  ( .A(\U1/aes_core/SB3/n1780 ), .B(
        \U1/aes_core/SB3/n1779 ), .Y(\U1/aes_core/SB3/n3297 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1394  ( .A(\U1/aes_core/SB3/n3297 ), .B(
        \U1/aes_core/SB3/n2021 ), .Y(\U1/aes_core/SB3/n1965 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1393  ( .A(\U1/aes_core/SB3/n3300 ), .B(
        \U1/aes_core/SB3/n2006 ), .Y(\U1/aes_core/SB3/n1878 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1392  ( .A(\U1/aes_core/SB3/n3333 ), .B(
        \U1/aes_core/SB3/n3305 ), .Y(\U1/aes_core/SB3/n1842 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1391  ( .A0(\U1/aes_core/SB3/n3300 ), 
        .A1(\U1/aes_core/SB3/n3342 ), .B0(\U1/aes_core/SB3/n1842 ), .Y(
        \U1/aes_core/SB3/n1787 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1390  ( .A(\U1/aes_core/SB3/n1912 ), .Y(
        \U1/aes_core/SB3/n3325 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1389  ( .A(\U1/aes_core/SB3/n3268 ), .B(
        \U1/aes_core/SB3/n3325 ), .Y(\U1/aes_core/SB3/n1977 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1388  ( .A(\U1/aes_core/SB3/n3268 ), .B(
        \U1/aes_core/SB3/n3334 ), .Y(\U1/aes_core/SB3/n1954 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1387  ( .A(\U1/aes_core/SB3/n1782 ), .B(
        \U1/aes_core/SB3/n1781 ), .Y(\U1/aes_core/SB3/n2008 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1386  ( .A(\U1/aes_core/SB3/n2008 ), .Y(
        \U1/aes_core/SB3/n3307 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1385  ( .A(\U1/aes_core/SB3/n3307 ), .B(
        \U1/aes_core/SB3/n2019 ), .Y(\U1/aes_core/SB3/n1855 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1384  ( .A(\U1/aes_core/SB3/n3307 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1902 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1383  ( .A(\U1/aes_core/SB3/n1977 ), .B(
        \U1/aes_core/SB3/n1954 ), .C(\U1/aes_core/SB3/n1855 ), .D(
        \U1/aes_core/SB3/n1902 ), .Y(\U1/aes_core/SB3/n1786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1382  ( .A(\U1/aes_core/SB3/n3346 ), .Y(
        \U1/aes_core/SB3/n3275 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1381  ( .A(\U1/aes_core/SB3/n3275 ), .B(
        \U1/aes_core/SB3/n1976 ), .Y(\U1/aes_core/SB3/n1927 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1380  ( .A(\U1/aes_core/SB3/n3297 ), .Y(
        \U1/aes_core/SB3/n3282 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1379  ( .A(\U1/aes_core/SB3/n1976 ), .B(
        \U1/aes_core/SB3/n3282 ), .Y(\U1/aes_core/SB3/n1922 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1378  ( .A(\U1/aes_core/SB3/n3322 ), .B(
        \U1/aes_core/SB3/n3276 ), .Y(\U1/aes_core/SB3/n1830 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1377  ( .A(\U1/aes_core/SB3/n3299 ), .B(
        \U1/aes_core/SB3/n2019 ), .Y(\U1/aes_core/SB3/n1909 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1376  ( .A(\U1/aes_core/SB3/n1927 ), .B(
        \U1/aes_core/SB3/n1922 ), .C(\U1/aes_core/SB3/n1830 ), .D(
        \U1/aes_core/SB3/n1909 ), .Y(\U1/aes_core/SB3/n1785 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1375  ( .A(\U1/aes_core/SB3/n3279 ), .Y(
        \U1/aes_core/SB3/n3323 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1374  ( .A(\U1/aes_core/SB3/n3274 ), .B(
        \U1/aes_core/SB3/n3323 ), .Y(\U1/aes_core/SB3/n1820 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1373  ( .A(\U1/aes_core/SB3/n2054 ), .B(
        \U1/aes_core/SB3/n3274 ), .Y(\U1/aes_core/SB3/n1864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1372  ( .A(\U1/aes_core/SB3/n1783 ), .B(
        \U1/aes_core/SB3/n1782 ), .Y(\U1/aes_core/SB3/n3303 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1371  ( .A(\U1/aes_core/SB3/n3303 ), .Y(
        \U1/aes_core/SB3/n3329 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1370  ( .A(\U1/aes_core/SB3/n2068 ), .B(
        \U1/aes_core/SB3/n3329 ), .Y(\U1/aes_core/SB3/n1890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1369  ( .A(\U1/aes_core/SB3/n2054 ), .B(
        \U1/aes_core/SB3/n3324 ), .Y(\U1/aes_core/SB3/n1990 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1368  ( .A(\U1/aes_core/SB3/n1820 ), .B(
        \U1/aes_core/SB3/n1864 ), .C(\U1/aes_core/SB3/n1890 ), .D(
        \U1/aes_core/SB3/n1990 ), .Y(\U1/aes_core/SB3/n1784 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1367  ( .A(\U1/aes_core/SB3/n1965 ), .B(
        \U1/aes_core/SB3/n1878 ), .C(\U1/aes_core/SB3/n1787 ), .D(
        \U1/aes_core/SB3/n1786 ), .E(\U1/aes_core/SB3/n1785 ), .F(
        \U1/aes_core/SB3/n1784 ), .Y(\U1/aes_core/SB3/n3286 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1366  ( .A(\U1/aes_core/SB3/n3279 ), .B(
        \U1/aes_core/SB3/n2021 ), .Y(\U1/aes_core/SB3/n1831 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1365  ( .A(\U1/aes_core/SB3/n3280 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n1980 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1364  ( .A(\U1/aes_core/SB3/n3278 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n1872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1363  ( .A(\U1/aes_core/SB3/n3278 ), .B(
        \U1/aes_core/SB3/n3281 ), .Y(\U1/aes_core/SB3/n1881 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1362  ( .A(\U1/aes_core/SB3/n3342 ), .B(
        \U1/aes_core/SB3/n3308 ), .Y(\U1/aes_core/SB3/n1919 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1361  ( .A(\U1/aes_core/SB3/n3307 ), .B(
        \U1/aes_core/SB3/n3325 ), .Y(\U1/aes_core/SB3/n1923 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1360  ( .A(\U1/aes_core/SB3/n2058 ), .B(
        \U1/aes_core/SB3/n3329 ), .Y(\U1/aes_core/SB3/n1844 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1359  ( .A(\U1/aes_core/SB3/n3331 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1857 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1358  ( .AN(\U1/aes_core/SB3/n1919 ), 
        .B(\U1/aes_core/SB3/n1923 ), .C(\U1/aes_core/SB3/n1844 ), .D(
        \U1/aes_core/SB3/n1857 ), .Y(\U1/aes_core/SB3/n1791 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1357  ( .A(\U1/aes_core/SB3/n3300 ), .B(
        \U1/aes_core/SB3/n3281 ), .Y(\U1/aes_core/SB3/n1891 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1356  ( .A(\U1/aes_core/SB3/n3347 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n1967 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1355  ( .A(\U1/aes_core/SB3/n1995 ), .B(
        \U1/aes_core/SB3/n3346 ), .Y(\U1/aes_core/SB3/n1930 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1354  ( .A(\U1/aes_core/SB3/n1995 ), .B(
        \U1/aes_core/SB3/n2006 ), .Y(\U1/aes_core/SB3/n1828 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1353  ( .A0(\U1/aes_core/SB3/n3281 ), 
        .A1(\U1/aes_core/SB3/n1995 ), .B0(\U1/aes_core/SB3/n3300 ), .B1(
        \U1/aes_core/SB3/n3346 ), .Y(\U1/aes_core/SB3/n1789 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1352  ( .A0(\U1/aes_core/SB3/n1888 ), 
        .A1(\U1/aes_core/SB3/n2070 ), .B0(\U1/aes_core/SB3/n2020 ), .B1(
        \U1/aes_core/SB3/n3280 ), .Y(\U1/aes_core/SB3/n1788 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1351  ( .A(\U1/aes_core/SB3/n1891 ), .B(
        \U1/aes_core/SB3/n1967 ), .C(\U1/aes_core/SB3/n1930 ), .D(
        \U1/aes_core/SB3/n1828 ), .E(\U1/aes_core/SB3/n1789 ), .F(
        \U1/aes_core/SB3/n1788 ), .Y(\U1/aes_core/SB3/n1790 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1350  ( .A(\U1/aes_core/SB3/n1831 ), .B(
        \U1/aes_core/SB3/n1980 ), .C(\U1/aes_core/SB3/n1872 ), .D(
        \U1/aes_core/SB3/n1881 ), .E(\U1/aes_core/SB3/n1791 ), .F(
        \U1/aes_core/SB3/n1790 ), .Y(\U1/aes_core/SB3/n3321 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U1349  ( .A1N(\U1/aes_core/SB3/n3299 ), 
        .A0(\U1/aes_core/SB3/n3343 ), .B0(\U1/aes_core/SB3/n2020 ), .Y(
        \U1/aes_core/SB3/n1792 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1348  ( .A(\U1/aes_core/SB3/n1995 ), .B(
        \U1/aes_core/SB3/n2039 ), .Y(\U1/aes_core/SB3/n1943 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1347  ( .A(\U1/aes_core/SB3/n3280 ), .B(
        \U1/aes_core/SB3/n2057 ), .Y(\U1/aes_core/SB3/n1850 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1346  ( .A(\U1/aes_core/SB3/n3280 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n1886 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1345  ( .A(\U1/aes_core/SB3/n1792 ), .B(
        \U1/aes_core/SB3/n1943 ), .C(\U1/aes_core/SB3/n1850 ), .D(
        \U1/aes_core/SB3/n1886 ), .Y(\U1/aes_core/SB3/n1797 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1344  ( .A0(\U1/aes_core/SB3/n2057 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n2021 ), .B1(
        \U1/aes_core/SB3/n3296 ), .C0(\U1/aes_core/SB3/n1912 ), .C1(
        \U1/aes_core/SB3/n3309 ), .Y(\U1/aes_core/SB3/n1796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1343  ( .A(\U1/aes_core/SB3/n3342 ), .B(
        \U1/aes_core/SB3/n3309 ), .Y(\U1/aes_core/SB3/n1972 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1342  ( .A(\U1/aes_core/SB3/n2065 ), .B(
        \U1/aes_core/SB3/n2010 ), .Y(\U1/aes_core/SB3/n1833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1341  ( .A(\U1/aes_core/SB3/n1833 ), .Y(
        \U1/aes_core/SB3/n1793 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1340  ( .A(\U1/aes_core/SB3/n3329 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1339  ( .A(\U1/aes_core/SB3/n1976 ), .B(
        \U1/aes_core/SB3/n2054 ), .Y(\U1/aes_core/SB3/n1853 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1338  ( .AN(\U1/aes_core/SB3/n1972 ), 
        .B(\U1/aes_core/SB3/n1793 ), .C(\U1/aes_core/SB3/n1866 ), .D(
        \U1/aes_core/SB3/n1853 ), .Y(\U1/aes_core/SB3/n1795 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1337  ( .A(\U1/aes_core/SB3/n1888 ), .B(
        \U1/aes_core/SB3/n2021 ), .Y(\U1/aes_core/SB3/n1918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1336  ( .A(\U1/aes_core/SB3/n1806 ), .B(
        \U1/aes_core/SB3/n3297 ), .Y(\U1/aes_core/SB3/n1895 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1335  ( .A(\U1/aes_core/SB3/n2008 ), .B(
        \U1/aes_core/SB3/n2020 ), .Y(\U1/aes_core/SB3/n1935 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1334  ( .A(\U1/aes_core/SB3/n2008 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n1827 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1333  ( .A(\U1/aes_core/SB3/n1918 ), .B(
        \U1/aes_core/SB3/n1895 ), .C(\U1/aes_core/SB3/n1935 ), .D(
        \U1/aes_core/SB3/n1827 ), .Y(\U1/aes_core/SB3/n1794 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1332  ( .A(\U1/aes_core/SB3/n1797 ), .B(
        \U1/aes_core/SB3/n1796 ), .C(\U1/aes_core/SB3/n1795 ), .D(
        \U1/aes_core/SB3/n1794 ), .Y(\U1/aes_core/SB3/n3293 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1331  ( .A(\U1/aes_core/SB3/n3308 ), .Y(
        \U1/aes_core/SB3/n3327 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1330  ( .A0(\U1/aes_core/SB3/n3330 ), 
        .A1(\U1/aes_core/SB3/n3268 ), .B0(\U1/aes_core/SB3/n2068 ), .B1(
        \U1/aes_core/SB3/n3327 ), .Y(\U1/aes_core/SB3/n1798 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1329  ( .A0(\U1/aes_core/SB3/n3297 ), 
        .A1(\U1/aes_core/SB3/n3347 ), .B0(\U1/aes_core/SB3/n3280 ), .B1(
        \U1/aes_core/SB3/n3346 ), .C0(\U1/aes_core/SB3/n1798 ), .Y(
        \U1/aes_core/SB3/n1804 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1328  ( .A(\U1/aes_core/SB3/n3303 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n1862 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1327  ( .A(\U1/aes_core/SB3/n3332 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1326  ( .A(\U1/aes_core/SB3/n3268 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1325  ( .A(\U1/aes_core/SB3/n3330 ), .B(
        \U1/aes_core/SB3/n3307 ), .Y(\U1/aes_core/SB3/n1839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1324  ( .AN(\U1/aes_core/SB3/n1862 ), 
        .B(\U1/aes_core/SB3/n1874 ), .C(\U1/aes_core/SB3/n1867 ), .D(
        \U1/aes_core/SB3/n1839 ), .Y(\U1/aes_core/SB3/n1803 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1323  ( .A(\U1/aes_core/SB3/n3281 ), .B(
        \U1/aes_core/SB3/n2057 ), .Y(\U1/aes_core/SB3/n1948 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1322  ( .A0(\U1/aes_core/SB3/n3325 ), 
        .A1(\U1/aes_core/SB3/n1948 ), .B0(\U1/aes_core/SB3/n3322 ), .Y(
        \U1/aes_core/SB3/n1801 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1321  ( .A(\U1/aes_core/SB3/n3344 ), .Y(
        \U1/aes_core/SB3/n1949 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1320  ( .A0(\U1/aes_core/SB3/n2058 ), 
        .A1(\U1/aes_core/SB3/n3323 ), .B0(\U1/aes_core/SB3/n1949 ), .Y(
        \U1/aes_core/SB3/n1800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1319  ( .A(\U1/aes_core/SB3/n2020 ), .Y(
        \U1/aes_core/SB3/n2060 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1318  ( .A0(\U1/aes_core/SB3/n1952 ), 
        .A1(\U1/aes_core/SB3/n1976 ), .B0(\U1/aes_core/SB3/n2060 ), .Y(
        \U1/aes_core/SB3/n1799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1317  ( .A(\U1/aes_core/SB3/n2058 ), .B(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n1925 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1316  ( .A(\U1/aes_core/SB3/n1801 ), .B(
        \U1/aes_core/SB3/n1800 ), .C(\U1/aes_core/SB3/n1799 ), .D(
        \U1/aes_core/SB3/n1925 ), .Y(\U1/aes_core/SB3/n1802 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1315  ( .A(\U1/aes_core/SB3/n3286 ), .B(
        \U1/aes_core/SB3/n3321 ), .C(\U1/aes_core/SB3/n3293 ), .D(
        \U1/aes_core/SB3/n1804 ), .E(\U1/aes_core/SB3/n1803 ), .F(
        \U1/aes_core/SB3/n1802 ), .Y(\U1/aes_core/SB3/n2074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1314  ( .A0(\U1/aes_core/SB3/n2019 ), 
        .A1(\U1/aes_core/SB3/n3330 ), .B0(\U1/aes_core/SB3/n3324 ), .Y(
        \U1/aes_core/SB3/n1805 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1313  ( .A(\U1/aes_core/SB3/n3269 ), .B(
        \U1/aes_core/SB3/n2058 ), .Y(\U1/aes_core/SB3/n1910 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1312  ( .A(\U1/aes_core/SB3/n2055 ), .B(
        \U1/aes_core/SB3/n3276 ), .Y(\U1/aes_core/SB3/n1819 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1311  ( .A(\U1/aes_core/SB3/n3340 ), .B(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n1921 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1310  ( .A(\U1/aes_core/SB3/n1805 ), .B(
        \U1/aes_core/SB3/n1910 ), .C(\U1/aes_core/SB3/n1819 ), .D(
        \U1/aes_core/SB3/n1921 ), .Y(\U1/aes_core/SB3/n1810 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1309  ( .A0(\U1/aes_core/SB3/n2020 ), 
        .A1(\U1/aes_core/SB3/n1806 ), .B0(\U1/aes_core/SB3/n3302 ), .B1(
        \U1/aes_core/SB3/n3347 ), .C0(\U1/aes_core/SB3/n3346 ), .C1(
        \U1/aes_core/SB3/n2065 ), .Y(\U1/aes_core/SB3/n1809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1308  ( .A(\U1/aes_core/SB3/n1976 ), .B(
        \U1/aes_core/SB3/n3334 ), .Y(\U1/aes_core/SB3/n1841 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1307  ( .A(\U1/aes_core/SB3/n2058 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1964 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1306  ( .A(\U1/aes_core/SB3/n3275 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1863 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1305  ( .A(\U1/aes_core/SB3/n3340 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1926 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1304  ( .A(\U1/aes_core/SB3/n1841 ), .B(
        \U1/aes_core/SB3/n1964 ), .C(\U1/aes_core/SB3/n1863 ), .D(
        \U1/aes_core/SB3/n1926 ), .Y(\U1/aes_core/SB3/n1808 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1303  ( .A(\U1/aes_core/SB3/n3340 ), .B(
        \U1/aes_core/SB3/n3332 ), .Y(\U1/aes_core/SB3/n1889 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1302  ( .A(\U1/aes_core/SB3/n3333 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n1876 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1301  ( .A(\U1/aes_core/SB3/n3274 ), .B(
        \U1/aes_core/SB3/n3276 ), .Y(\U1/aes_core/SB3/n1854 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1300  ( .A(\U1/aes_core/SB3/n3323 ), .B(
        \U1/aes_core/SB3/n3327 ), .Y(\U1/aes_core/SB3/n1829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1299  ( .A(\U1/aes_core/SB3/n1889 ), .B(
        \U1/aes_core/SB3/n1876 ), .C(\U1/aes_core/SB3/n1854 ), .D(
        \U1/aes_core/SB3/n1829 ), .Y(\U1/aes_core/SB3/n1807 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1298  ( .A(\U1/aes_core/SB3/n1810 ), .B(
        \U1/aes_core/SB3/n1809 ), .C(\U1/aes_core/SB3/n1808 ), .D(
        \U1/aes_core/SB3/n1807 ), .Y(\U1/aes_core/SB3/n1811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1297  ( .A(\U1/aes_core/SB3/n1811 ), .Y(
        \U1/aes_core/SB3/n3284 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1296  ( .A0(\U1/aes_core/SB3/n3308 ), 
        .A1(\U1/aes_core/SB3/n2039 ), .B0(\U1/aes_core/SB3/n3297 ), .B1(
        \U1/aes_core/SB3/n2070 ), .C0(\U1/aes_core/SB3/n3284 ), .Y(
        \U1/aes_core/SB3/n1818 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1295  ( .A(\U1/aes_core/SB3/n3329 ), .B(
        \U1/aes_core/SB3/n3274 ), .Y(\U1/aes_core/SB3/n1920 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U1294  ( .A1N(\U1/aes_core/SB3/n1920 ), 
        .A0(\U1/aes_core/SB3/n3305 ), .B0(\U1/aes_core/SB3/n2019 ), .Y(
        \U1/aes_core/SB3/n1814 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1293  ( .A(\U1/aes_core/SB3/n2017 ), .B(
        \U1/aes_core/SB3/n3346 ), .Y(\U1/aes_core/SB3/n2018 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1292  ( .A0(\U1/aes_core/SB3/n3331 ), 
        .A1(\U1/aes_core/SB3/n2018 ), .B0(\U1/aes_core/SB3/n3268 ), .Y(
        \U1/aes_core/SB3/n1813 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1291  ( .A0(\U1/aes_core/SB3/n2058 ), 
        .A1(\U1/aes_core/SB3/n3333 ), .B0(\U1/aes_core/SB3/n2055 ), .Y(
        \U1/aes_core/SB3/n1812 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1290  ( .A(\U1/aes_core/SB3/n2054 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n1851 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1289  ( .A(\U1/aes_core/SB3/n1814 ), .B(
        \U1/aes_core/SB3/n1813 ), .C(\U1/aes_core/SB3/n1812 ), .D(
        \U1/aes_core/SB3/n1851 ), .Y(\U1/aes_core/SB3/n1817 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1288  ( .A(\U1/aes_core/SB3/n3275 ), .B(
        \U1/aes_core/SB3/n2060 ), .Y(\U1/aes_core/SB3/n2059 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1287  ( .A(\U1/aes_core/SB3/n2053 ), .B(
        \U1/aes_core/SB3/n1976 ), .Y(\U1/aes_core/SB3/n1815 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1286  ( .A0(\U1/aes_core/SB3/n2059 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n1815 ), .B1(
        \U1/aes_core/SB3/n2010 ), .C0(\U1/aes_core/SB3/n3302 ), .C1(
        \U1/aes_core/SB3/n3278 ), .Y(\U1/aes_core/SB3/n1816 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1285  ( .A(\U1/aes_core/SB3/n3353 ), .B(
        \U1/aes_core/SB3/n3295 ), .C(\U1/aes_core/SB3/n2074 ), .D(
        \U1/aes_core/SB3/n1818 ), .E(\U1/aes_core/SB3/n1817 ), .F(
        \U1/aes_core/SB3/n1816 ), .Y(\U1/aes_core/sb3 [10]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1284  ( .A(\U1/aes_core/SB3/n3347 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n2034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1283  ( .A(\U1/aes_core/SB3/n3330 ), .B(
        \U1/aes_core/SB3/n1952 ), .Y(\U1/aes_core/SB3/n2036 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1282  ( .AN(\U1/aes_core/SB3/n1821 ), 
        .B(\U1/aes_core/SB3/n1820 ), .C(\U1/aes_core/SB3/n1819 ), .D(
        \U1/aes_core/SB3/n2036 ), .Y(\U1/aes_core/SB3/n1826 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1281  ( .A(\U1/aes_core/SB3/n3324 ), .B(
        \U1/aes_core/SB3/n2055 ), .Y(\U1/aes_core/SB3/n1983 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1280  ( .A0(\U1/aes_core/SB3/n3269 ), 
        .A1(\U1/aes_core/SB3/n3268 ), .B0(\U1/aes_core/SB3/n3323 ), .Y(
        \U1/aes_core/SB3/n1822 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1279  ( .A(\U1/aes_core/SB3/n3340 ), .B(
        \U1/aes_core/SB3/n1952 ), .Y(\U1/aes_core/SB3/n2061 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U1278  ( .A0(\U1/aes_core/SB3/n1983 ), 
        .A1(\U1/aes_core/SB3/n3296 ), .B0(\U1/aes_core/SB3/n1822 ), .C0(
        \U1/aes_core/SB3/n2061 ), .Y(\U1/aes_core/SB3/n1825 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1277  ( .A0(\U1/aes_core/SB3/n2020 ), 
        .A1(\U1/aes_core/SB3/n2070 ), .B0(\U1/aes_core/SB3/n1823 ), .B1(
        \U1/aes_core/SB3/n3308 ), .C0(\U1/aes_core/SB3/n3281 ), .C1(
        \U1/aes_core/SB3/n2065 ), .Y(\U1/aes_core/SB3/n1824 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1276  ( .A(\U1/aes_core/SB3/n1828 ), .B(
        \U1/aes_core/SB3/n2034 ), .C(\U1/aes_core/SB3/n1827 ), .D(
        \U1/aes_core/SB3/n1826 ), .E(\U1/aes_core/SB3/n1825 ), .F(
        \U1/aes_core/SB3/n1824 ), .Y(\U1/aes_core/SB3/n1962 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1275  ( .A(\U1/aes_core/SB3/n3323 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n2040 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1274  ( .AN(\U1/aes_core/SB3/n1831 ), 
        .B(\U1/aes_core/SB3/n1830 ), .C(\U1/aes_core/SB3/n1829 ), .D(
        \U1/aes_core/SB3/n2040 ), .Y(\U1/aes_core/SB3/n1838 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U1273  ( .A0(\U1/aes_core/SB3/n3331 ), 
        .A1(\U1/aes_core/SB3/n3327 ), .B0(\U1/aes_core/SB3/n3332 ), .B1(
        \U1/aes_core/SB3/n3334 ), .C0(\U1/aes_core/SB3/n3274 ), .C1(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n1837 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1272  ( .A0(\U1/aes_core/SB3/n3301 ), 
        .A1(\U1/aes_core/SB3/n3280 ), .B0(\U1/aes_core/SB3/n2021 ), .B1(
        \U1/aes_core/SB3/n2020 ), .Y(\U1/aes_core/SB3/n1832 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1271  ( .A0(\U1/aes_core/SB3/n1952 ), 
        .A1(\U1/aes_core/SB3/n3323 ), .B0(\U1/aes_core/SB3/n3276 ), .B1(
        \U1/aes_core/SB3/n3299 ), .C0(\U1/aes_core/SB3/n1832 ), .Y(
        \U1/aes_core/SB3/n1836 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1270  ( .A(\U1/aes_core/SB3/n3308 ), .B(
        \U1/aes_core/SB3/n3343 ), .Y(\U1/aes_core/SB3/n3270 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1269  ( .A(\U1/aes_core/SB3/n3344 ), .B(
        \U1/aes_core/SB3/n3347 ), .Y(\U1/aes_core/SB3/n1834 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1268  ( .A0(\U1/aes_core/SB3/n3340 ), 
        .A1(\U1/aes_core/SB3/n3270 ), .B0(\U1/aes_core/SB3/n2058 ), .B1(
        \U1/aes_core/SB3/n1834 ), .C0(\U1/aes_core/SB3/n1833 ), .Y(
        \U1/aes_core/SB3/n1835 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1267  ( .AN(\U1/aes_core/SB3/n1838 ), 
        .B(\U1/aes_core/SB3/n1837 ), .C(\U1/aes_core/SB3/n1836 ), .D(
        \U1/aes_core/SB3/n1835 ), .Y(\U1/aes_core/SB3/n1988 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1266  ( .A(\U1/aes_core/SB3/n1995 ), .B(
        \U1/aes_core/SB3/n3302 ), .Y(\U1/aes_core/SB3/n2024 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1265  ( .A0(\U1/aes_core/SB3/n3303 ), 
        .A1(\U1/aes_core/SB3/n3302 ), .B0(\U1/aes_core/SB3/n1839 ), .Y(
        \U1/aes_core/SB3/n1849 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1264  ( .A0(\U1/aes_core/SB3/n2058 ), 
        .A1(\U1/aes_core/SB3/n3332 ), .B0(\U1/aes_core/SB3/n3275 ), .B1(
        \U1/aes_core/SB3/n3307 ), .Y(\U1/aes_core/SB3/n1840 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1263  ( .A0(\U1/aes_core/SB3/n3344 ), 
        .A1(\U1/aes_core/SB3/n2039 ), .B0(\U1/aes_core/SB3/n2057 ), .B1(
        \U1/aes_core/SB3/n3343 ), .C0(\U1/aes_core/SB3/n1840 ), .Y(
        \U1/aes_core/SB3/n1848 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1262  ( .A(\U1/aes_core/SB3/n1912 ), .B(
        \U1/aes_core/SB3/n3308 ), .Y(\U1/aes_core/SB3/n3292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1261  ( .A(\U1/aes_core/SB3/n3305 ), .B(
        \U1/aes_core/SB3/n3323 ), .Y(\U1/aes_core/SB3/n2037 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1260  ( .AN(\U1/aes_core/SB3/n3292 ), 
        .B(\U1/aes_core/SB3/n1842 ), .C(\U1/aes_core/SB3/n1841 ), .D(
        \U1/aes_core/SB3/n2037 ), .Y(\U1/aes_core/SB3/n1847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1259  ( .A(\U1/aes_core/SB3/n3280 ), .B(
        \U1/aes_core/SB3/n3297 ), .Y(\U1/aes_core/SB3/n2015 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1258  ( .AN(\U1/aes_core/SB3/n2015 ), 
        .B(\U1/aes_core/SB3/n1845 ), .C(\U1/aes_core/SB3/n1844 ), .D(
        \U1/aes_core/SB3/n1843 ), .Y(\U1/aes_core/SB3/n1846 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1257  ( .A(\U1/aes_core/SB3/n2024 ), .B(
        \U1/aes_core/SB3/n1850 ), .C(\U1/aes_core/SB3/n1849 ), .D(
        \U1/aes_core/SB3/n1848 ), .E(\U1/aes_core/SB3/n1847 ), .F(
        \U1/aes_core/SB3/n1846 ), .Y(\U1/aes_core/SB3/n1924 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1256  ( .A(\U1/aes_core/SB3/n2017 ), .B(
        \U1/aes_core/SB3/n3300 ), .Y(\U1/aes_core/SB3/n2064 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1255  ( .A0(\U1/aes_core/SB3/n2017 ), 
        .A1(\U1/aes_core/SB3/n3280 ), .B0(\U1/aes_core/SB3/n1851 ), .Y(
        \U1/aes_core/SB3/n1861 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1254  ( .A(\U1/aes_core/SB3/n3343 ), .B(
        \U1/aes_core/SB3/n1912 ), .Y(\U1/aes_core/SB3/n2023 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1253  ( .A(\U1/aes_core/SB3/n1949 ), .B(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n3312 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1252  ( .AN(\U1/aes_core/SB3/n2023 ), 
        .B(\U1/aes_core/SB3/n1853 ), .C(\U1/aes_core/SB3/n1852 ), .D(
        \U1/aes_core/SB3/n3312 ), .Y(\U1/aes_core/SB3/n1860 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1251  ( .A(\U1/aes_core/SB3/n3274 ), .B(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n2045 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1250  ( .A(\U1/aes_core/SB3/n3339 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n3267 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1249  ( .A(\U1/aes_core/SB3/n2019 ), .B(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n3335 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1248  ( .A(\U1/aes_core/SB3/n1854 ), .B(
        \U1/aes_core/SB3/n2045 ), .C(\U1/aes_core/SB3/n3267 ), .D(
        \U1/aes_core/SB3/n3335 ), .Y(\U1/aes_core/SB3/n1859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1247  ( .A(\U1/aes_core/SB3/n3322 ), .B(
        \U1/aes_core/SB3/n3333 ), .Y(\U1/aes_core/SB3/n2005 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1246  ( .A(\U1/aes_core/SB3/n1857 ), .B(
        \U1/aes_core/SB3/n1856 ), .C(\U1/aes_core/SB3/n2005 ), .D(
        \U1/aes_core/SB3/n1855 ), .Y(\U1/aes_core/SB3/n1858 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1245  ( .A(\U1/aes_core/SB3/n2064 ), .B(
        \U1/aes_core/SB3/n1862 ), .C(\U1/aes_core/SB3/n1861 ), .D(
        \U1/aes_core/SB3/n1860 ), .E(\U1/aes_core/SB3/n1859 ), .F(
        \U1/aes_core/SB3/n1858 ), .Y(\U1/aes_core/SB3/n1940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1244  ( .A(\U1/aes_core/SB3/n3302 ), .B(
        \U1/aes_core/SB3/n2021 ), .Y(\U1/aes_core/SB3/n2016 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1243  ( .A(\U1/aes_core/SB3/n3324 ), .B(
        \U1/aes_core/SB3/n3331 ), .Y(\U1/aes_core/SB3/n2041 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1242  ( .A(\U1/aes_core/SB3/n3334 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n3265 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1241  ( .A(\U1/aes_core/SB3/n1864 ), .B(
        \U1/aes_core/SB3/n1863 ), .C(\U1/aes_core/SB3/n2041 ), .D(
        \U1/aes_core/SB3/n3265 ), .Y(\U1/aes_core/SB3/n1871 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1240  ( .A(\U1/aes_core/SB3/n1952 ), .B(
        \U1/aes_core/SB3/n3276 ), .Y(\U1/aes_core/SB3/n2027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1239  ( .A(\U1/aes_core/SB3/n3333 ), .B(
        \U1/aes_core/SB3/n1952 ), .Y(\U1/aes_core/SB3/n3311 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1238  ( .A(\U1/aes_core/SB3/n1866 ), .B(
        \U1/aes_core/SB3/n2027 ), .C(\U1/aes_core/SB3/n1865 ), .D(
        \U1/aes_core/SB3/n3311 ), .Y(\U1/aes_core/SB3/n1870 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U1237  ( .A(\U1/aes_core/SB3/n2055 ), .B(
        \U1/aes_core/SB3/n3329 ), .C(\U1/aes_core/SB3/n2053 ), .Y(
        \U1/aes_core/SB3/n1868 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1236  ( .A0(\U1/aes_core/SB3/n1868 ), 
        .A1(\U1/aes_core/SB3/n2010 ), .B0(\U1/aes_core/SB3/n2020 ), .B1(
        \U1/aes_core/SB3/n3347 ), .C0(\U1/aes_core/SB3/n1867 ), .Y(
        \U1/aes_core/SB3/n1869 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1235  ( .A(\U1/aes_core/SB3/n2016 ), .B(
        \U1/aes_core/SB3/n1873 ), .C(\U1/aes_core/SB3/n1872 ), .D(
        \U1/aes_core/SB3/n1871 ), .E(\U1/aes_core/SB3/n1870 ), .F(
        \U1/aes_core/SB3/n1869 ), .Y(\U1/aes_core/SB3/n1973 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1234  ( .A(\U1/aes_core/SB3/n3300 ), .B(
        \U1/aes_core/SB3/n1888 ), .Y(\U1/aes_core/SB3/n2028 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1233  ( .A0(\U1/aes_core/SB3/n2020 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n1874 ), .Y(
        \U1/aes_core/SB3/n1885 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1232  ( .A0(\U1/aes_core/SB3/n1976 ), 
        .A1(\U1/aes_core/SB3/n2019 ), .B0(\U1/aes_core/SB3/n3322 ), .B1(
        \U1/aes_core/SB3/n3334 ), .Y(\U1/aes_core/SB3/n1875 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1231  ( .A0(\U1/aes_core/SB3/n3308 ), 
        .A1(\U1/aes_core/SB3/n3346 ), .B0(\U1/aes_core/SB3/n3303 ), .B1(
        \U1/aes_core/SB3/n3279 ), .C0(\U1/aes_core/SB3/n1875 ), .Y(
        \U1/aes_core/SB3/n1884 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1230  ( .A(\U1/aes_core/SB3/n3303 ), .B(
        \U1/aes_core/SB3/n2020 ), .Y(\U1/aes_core/SB3/n3291 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1229  ( .A(\U1/aes_core/SB3/n3291 ), .Y(
        \U1/aes_core/SB3/n1877 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1228  ( .A(\U1/aes_core/SB3/n3332 ), .B(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n2047 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1227  ( .AN(\U1/aes_core/SB3/n1878 ), 
        .B(\U1/aes_core/SB3/n1877 ), .C(\U1/aes_core/SB3/n1876 ), .D(
        \U1/aes_core/SB3/n2047 ), .Y(\U1/aes_core/SB3/n1883 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1226  ( .A(\U1/aes_core/SB3/n2058 ), .B(
        \U1/aes_core/SB3/n3307 ), .Y(\U1/aes_core/SB3/n2003 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1225  ( .AN(\U1/aes_core/SB3/n1881 ), 
        .B(\U1/aes_core/SB3/n1880 ), .C(\U1/aes_core/SB3/n1879 ), .D(
        \U1/aes_core/SB3/n2003 ), .Y(\U1/aes_core/SB3/n1882 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1224  ( .A(\U1/aes_core/SB3/n2028 ), .B(
        \U1/aes_core/SB3/n1886 ), .C(\U1/aes_core/SB3/n1885 ), .D(
        \U1/aes_core/SB3/n1884 ), .E(\U1/aes_core/SB3/n1883 ), .F(
        \U1/aes_core/SB3/n1882 ), .Y(\U1/aes_core/SB3/n1947 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1223  ( .A0(\U1/aes_core/SB3/n2053 ), 
        .A1(\U1/aes_core/SB3/n2018 ), .B0(\U1/aes_core/SB3/n1976 ), .B1(
        \U1/aes_core/SB3/n2060 ), .Y(\U1/aes_core/SB3/n1887 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1222  ( .A0(\U1/aes_core/SB3/n3281 ), 
        .A1(\U1/aes_core/SB3/n3280 ), .B0(\U1/aes_core/SB3/n1888 ), .B1(
        \U1/aes_core/SB3/n3343 ), .C0(\U1/aes_core/SB3/n1887 ), .Y(
        \U1/aes_core/SB3/n1898 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1221  ( .A(\U1/aes_core/SB3/n3329 ), .B(
        \U1/aes_core/SB3/n3325 ), .Y(\U1/aes_core/SB3/n2044 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1220  ( .AN(\U1/aes_core/SB3/n1891 ), 
        .B(\U1/aes_core/SB3/n1890 ), .C(\U1/aes_core/SB3/n1889 ), .D(
        \U1/aes_core/SB3/n2044 ), .Y(\U1/aes_core/SB3/n1897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1219  ( .A0(\U1/aes_core/SB3/n3282 ), 
        .A1(\U1/aes_core/SB3/n3340 ), .B0(\U1/aes_core/SB3/n3322 ), .Y(
        \U1/aes_core/SB3/n1894 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1218  ( .A(\U1/aes_core/SB3/n3344 ), .B(
        \U1/aes_core/SB3/n1995 ), .Y(\U1/aes_core/SB3/n1892 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1217  ( .A0(\U1/aes_core/SB3/n3333 ), 
        .A1(\U1/aes_core/SB3/n1892 ), .B0(\U1/aes_core/SB3/n3329 ), .B1(
        \U1/aes_core/SB3/n1948 ), .Y(\U1/aes_core/SB3/n1893 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1216  ( .AN(\U1/aes_core/SB3/n1895 ), 
        .B(\U1/aes_core/SB3/n1894 ), .C(\U1/aes_core/SB3/n1893 ), .Y(
        \U1/aes_core/SB3/n1896 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1215  ( .A(\U1/aes_core/SB3/n1940 ), .B(
        \U1/aes_core/SB3/n1973 ), .C(\U1/aes_core/SB3/n1947 ), .D(
        \U1/aes_core/SB3/n1898 ), .E(\U1/aes_core/SB3/n1897 ), .F(
        \U1/aes_core/SB3/n1896 ), .Y(\U1/aes_core/SB3/n1999 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1214  ( .A(\U1/aes_core/SB3/n1962 ), .B(
        \U1/aes_core/SB3/n1988 ), .C(\U1/aes_core/SB3/n1924 ), .D(
        \U1/aes_core/SB3/n1999 ), .Y(\U1/aes_core/SB3/n1908 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1213  ( .A(\U1/aes_core/SB3/n3333 ), .B(
        \U1/aes_core/SB3/n2068 ), .Y(\U1/aes_core/SB3/n2009 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1212  ( .A(\U1/aes_core/SB3/n3323 ), .B(
        \U1/aes_core/SB3/n2060 ), .Y(\U1/aes_core/SB3/n2002 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1211  ( .A(\U1/aes_core/SB3/n3297 ), .B(
        \U1/aes_core/SB3/n3302 ), .Y(\U1/aes_core/SB3/n3306 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1210  ( .A0(\U1/aes_core/SB3/n1952 ), 
        .A1(\U1/aes_core/SB3/n3275 ), .B0(\U1/aes_core/SB3/n3306 ), .B1(
        \U1/aes_core/SB3/n3305 ), .Y(\U1/aes_core/SB3/n1899 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1209  ( .A0(\U1/aes_core/SB3/n2021 ), 
        .A1(\U1/aes_core/SB3/n2009 ), .B0(\U1/aes_core/SB3/n3278 ), .B1(
        \U1/aes_core/SB3/n2002 ), .C0(\U1/aes_core/SB3/n1899 ), .Y(
        \U1/aes_core/SB3/n1900 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1208  ( .A(\U1/aes_core/SB3/n1900 ), .Y(
        \U1/aes_core/SB3/n1907 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1207  ( .A0(\U1/aes_core/SB3/n3301 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n2020 ), .B1(
        \U1/aes_core/SB3/n1995 ), .Y(\U1/aes_core/SB3/n1901 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1206  ( .A0(\U1/aes_core/SB3/n2054 ), 
        .A1(\U1/aes_core/SB3/n3268 ), .B0(\U1/aes_core/SB3/n3327 ), .B1(
        \U1/aes_core/SB3/n3282 ), .C0(\U1/aes_core/SB3/n1901 ), .Y(
        \U1/aes_core/SB3/n1906 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1205  ( .A0(\U1/aes_core/SB3/n2068 ), 
        .A1(\U1/aes_core/SB3/n3323 ), .B0(\U1/aes_core/SB3/n2055 ), .Y(
        \U1/aes_core/SB3/n1904 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1204  ( .A(\U1/aes_core/SB3/n3340 ), .B(
        \U1/aes_core/SB3/n3305 ), .Y(\U1/aes_core/SB3/n2026 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB3/U1203  ( .A(\U1/aes_core/SB3/n1904 ), .B(
        \U1/aes_core/SB3/n2026 ), .C(\U1/aes_core/SB3/n1903 ), .D(
        \U1/aes_core/SB3/n1902 ), .Y(\U1/aes_core/SB3/n1905 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1202  ( .AN(\U1/aes_core/SB3/n1908 ), 
        .B(\U1/aes_core/SB3/n1907 ), .C(\U1/aes_core/SB3/n1906 ), .D(
        \U1/aes_core/SB3/n1905 ), .Y(\U1/aes_core/sb3 [11]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1201  ( .A0(\U1/aes_core/SB3/n1920 ), 
        .A1(\U1/aes_core/SB3/n2008 ), .B0(\U1/aes_core/SB3/n3297 ), .Y(
        \U1/aes_core/SB3/n1917 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1200  ( .A(\U1/aes_core/SB3/n1949 ), .B(
        \U1/aes_core/SB3/n3325 ), .Y(\U1/aes_core/SB3/n2035 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U1199  ( .A(\U1/aes_core/SB3/n1910 ), .B(
        \U1/aes_core/SB3/n2035 ), .C(\U1/aes_core/SB3/n1909 ), .Y(
        \U1/aes_core/SB3/n1916 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1198  ( .A(\U1/aes_core/SB3/n2053 ), .B(
        \U1/aes_core/SB3/n3322 ), .Y(\U1/aes_core/SB3/n1913 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1197  ( .A(\U1/aes_core/SB3/n3305 ), .B(
        \U1/aes_core/SB3/n1952 ), .Y(\U1/aes_core/SB3/n1911 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1196  ( .A0(\U1/aes_core/SB3/n1913 ), 
        .A1(\U1/aes_core/SB3/n1912 ), .B0(\U1/aes_core/SB3/n1911 ), .B1(
        \U1/aes_core/SB3/n2057 ), .C0(\U1/aes_core/SB3/n2006 ), .C1(
        \U1/aes_core/SB3/n2008 ), .Y(\U1/aes_core/SB3/n1915 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1195  ( .A0(\U1/aes_core/SB3/n3303 ), 
        .A1(\U1/aes_core/SB3/n2017 ), .B0(\U1/aes_core/SB3/n3281 ), .B1(
        \U1/aes_core/SB3/n3343 ), .C0(\U1/aes_core/SB3/n3308 ), .C1(
        \U1/aes_core/SB3/n2010 ), .Y(\U1/aes_core/SB3/n1914 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1194  ( .A(\U1/aes_core/SB3/n1919 ), .B(
        \U1/aes_core/SB3/n1918 ), .C(\U1/aes_core/SB3/n1917 ), .D(
        \U1/aes_core/SB3/n1916 ), .E(\U1/aes_core/SB3/n1915 ), .F(
        \U1/aes_core/SB3/n1914 ), .Y(\U1/aes_core/SB3/n2000 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1193  ( .A0(\U1/aes_core/SB3/n1920 ), 
        .A1(\U1/aes_core/SB3/n3280 ), .B0(\U1/aes_core/SB3/n3346 ), .Y(
        \U1/aes_core/SB3/n1946 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB3/U1192  ( .A0(\U1/aes_core/SB3/n3296 ), 
        .A1(\U1/aes_core/SB3/n3279 ), .A2(\U1/aes_core/SB3/n2010 ), .B0(
        \U1/aes_core/SB3/n3309 ), .Y(\U1/aes_core/SB3/n1945 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1191  ( .A(\U1/aes_core/SB3/n3276 ), .B(
        \U1/aes_core/SB3/n3327 ), .Y(\U1/aes_core/SB3/n2042 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1190  ( .A(\U1/aes_core/SB3/n1923 ), .B(
        \U1/aes_core/SB3/n1922 ), .C(\U1/aes_core/SB3/n1921 ), .D(
        \U1/aes_core/SB3/n2042 ), .Y(\U1/aes_core/SB3/n1942 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1189  ( .A(\U1/aes_core/SB3/n1924 ), .Y(
        \U1/aes_core/SB3/n1939 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1188  ( .A(\U1/aes_core/SB3/n3309 ), .B(
        \U1/aes_core/SB3/n3302 ), .Y(\U1/aes_core/SB3/n2022 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1187  ( .A0(\U1/aes_core/SB3/n2002 ), 
        .A1(\U1/aes_core/SB3/n2065 ), .B0(\U1/aes_core/SB3/n1925 ), .Y(
        \U1/aes_core/SB3/n1934 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1186  ( .A0(\U1/aes_core/SB3/n3280 ), 
        .A1(\U1/aes_core/SB3/n3342 ), .B0(\U1/aes_core/SB3/n3297 ), .B1(
        \U1/aes_core/SB3/n1995 ), .C0(\U1/aes_core/SB3/n3281 ), .C1(
        \U1/aes_core/SB3/n3309 ), .Y(\U1/aes_core/SB3/n1933 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1185  ( .A(\U1/aes_core/SB3/n3307 ), .B(
        \U1/aes_core/SB3/n3323 ), .Y(\U1/aes_core/SB3/n2046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1184  ( .A(\U1/aes_core/SB3/n2068 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n3272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1183  ( .A(\U1/aes_core/SB3/n1927 ), .B(
        \U1/aes_core/SB3/n1926 ), .C(\U1/aes_core/SB3/n2046 ), .D(
        \U1/aes_core/SB3/n3272 ), .Y(\U1/aes_core/SB3/n1932 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1182  ( .A(\U1/aes_core/SB3/n3333 ), .B(
        \U1/aes_core/SB3/n3299 ), .Y(\U1/aes_core/SB3/n2004 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1181  ( .AN(\U1/aes_core/SB3/n1930 ), 
        .B(\U1/aes_core/SB3/n1929 ), .C(\U1/aes_core/SB3/n1928 ), .D(
        \U1/aes_core/SB3/n2004 ), .Y(\U1/aes_core/SB3/n1931 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1180  ( .A(\U1/aes_core/SB3/n2022 ), .B(
        \U1/aes_core/SB3/n1935 ), .C(\U1/aes_core/SB3/n1934 ), .D(
        \U1/aes_core/SB3/n1933 ), .E(\U1/aes_core/SB3/n1932 ), .F(
        \U1/aes_core/SB3/n1931 ), .Y(\U1/aes_core/SB3/n1936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1179  ( .A(\U1/aes_core/SB3/n1936 ), .Y(
        \U1/aes_core/SB3/n1989 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1178  ( .A0(\U1/aes_core/SB3/n3344 ), 
        .A1(\U1/aes_core/SB3/n2017 ), .B0(\U1/aes_core/SB3/n3281 ), .B1(
        \U1/aes_core/SB3/n3347 ), .Y(\U1/aes_core/SB3/n1937 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U1177  ( .A0(\U1/aes_core/SB3/n3324 ), 
        .A1(\U1/aes_core/SB3/n3323 ), .B0(\U1/aes_core/SB3/n3330 ), .B1(
        \U1/aes_core/SB3/n3299 ), .C0(\U1/aes_core/SB3/n1937 ), .Y(
        \U1/aes_core/SB3/n1938 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1176  ( .AN(\U1/aes_core/SB3/n1940 ), 
        .B(\U1/aes_core/SB3/n1939 ), .C(\U1/aes_core/SB3/n1989 ), .D(
        \U1/aes_core/SB3/n1938 ), .Y(\U1/aes_core/SB3/n1941 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1175  ( .A(\U1/aes_core/SB3/n1946 ), .B(
        \U1/aes_core/SB3/n1945 ), .C(\U1/aes_core/SB3/n1944 ), .D(
        \U1/aes_core/SB3/n1943 ), .E(\U1/aes_core/SB3/n1942 ), .F(
        \U1/aes_core/SB3/n1941 ), .Y(\U1/aes_core/SB3/n1987 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1174  ( .A(\U1/aes_core/SB3/n1947 ), .Y(
        \U1/aes_core/SB3/n1951 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1173  ( .A0(\U1/aes_core/SB3/n1949 ), 
        .A1(\U1/aes_core/SB3/n1948 ), .B0(\U1/aes_core/SB3/n1952 ), .B1(
        \U1/aes_core/SB3/n3339 ), .Y(\U1/aes_core/SB3/n1950 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U1172  ( .A0(\U1/aes_core/SB3/n2006 ), 
        .A1(\U1/aes_core/SB3/n3309 ), .B0(\U1/aes_core/SB3/n1951 ), .C0(
        \U1/aes_core/SB3/n1950 ), .Y(\U1/aes_core/SB3/n1961 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1171  ( .A0(\U1/aes_core/SB3/n3276 ), 
        .A1(\U1/aes_core/SB3/n3275 ), .B0(\U1/aes_core/SB3/n3332 ), .Y(
        \U1/aes_core/SB3/n1956 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1170  ( .A0(\U1/aes_core/SB3/n1952 ), 
        .A1(\U1/aes_core/SB3/n3268 ), .B0(\U1/aes_core/SB3/n2060 ), .Y(
        \U1/aes_core/SB3/n1955 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1169  ( .A(\U1/aes_core/SB3/n1956 ), .B(
        \U1/aes_core/SB3/n1955 ), .C(\U1/aes_core/SB3/n1954 ), .D(
        \U1/aes_core/SB3/n1953 ), .Y(\U1/aes_core/SB3/n1960 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1168  ( .A(\U1/aes_core/SB3/n3325 ), .B(
        \U1/aes_core/SB3/n3334 ), .Y(\U1/aes_core/SB3/n1958 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1167  ( .A(\U1/aes_core/SB3/n3331 ), .B(
        \U1/aes_core/SB3/n3333 ), .Y(\U1/aes_core/SB3/n1957 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1166  ( .A(\U1/aes_core/SB3/n1976 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n3310 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1165  ( .A0(\U1/aes_core/SB3/n1958 ), 
        .A1(\U1/aes_core/SB3/n2070 ), .B0(\U1/aes_core/SB3/n1957 ), .B1(
        \U1/aes_core/SB3/n2008 ), .C0(\U1/aes_core/SB3/n3310 ), .C1(
        \U1/aes_core/SB3/n2039 ), .Y(\U1/aes_core/SB3/n1959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1164  ( .A(\U1/aes_core/SB3/n2000 ), .B(
        \U1/aes_core/SB3/n1987 ), .C(\U1/aes_core/SB3/n1962 ), .D(
        \U1/aes_core/SB3/n1961 ), .E(\U1/aes_core/SB3/n1960 ), .F(
        \U1/aes_core/SB3/n1959 ), .Y(\U1/aes_core/sb3 [12]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1163  ( .A(\U1/aes_core/SB3/n3300 ), .B(
        \U1/aes_core/SB3/n3297 ), .Y(\U1/aes_core/SB3/n2025 ) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U1162  ( .A1N(\U1/aes_core/SB3/n3306 ), 
        .A0(\U1/aes_core/SB3/n3279 ), .B0(\U1/aes_core/SB3/n3344 ), .Y(
        \U1/aes_core/SB3/n1971 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1161  ( .A(\U1/aes_core/SB3/n2053 ), .B(
        \U1/aes_core/SB3/n3268 ), .Y(\U1/aes_core/SB3/n1963 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1160  ( .A0(\U1/aes_core/SB3/n2070 ), 
        .A1(\U1/aes_core/SB3/n3302 ), .B0(\U1/aes_core/SB3/n1963 ), .B1(
        \U1/aes_core/SB3/n3281 ), .C0(\U1/aes_core/SB3/n3297 ), .C1(
        \U1/aes_core/SB3/n3278 ), .Y(\U1/aes_core/SB3/n1970 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1159  ( .A(\U1/aes_core/SB3/n3327 ), .B(
        \U1/aes_core/SB3/n2019 ), .Y(\U1/aes_core/SB3/n2043 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1158  ( .A(\U1/aes_core/SB3/n3299 ), .B(
        \U1/aes_core/SB3/n3282 ), .Y(\U1/aes_core/SB3/n3266 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1157  ( .AN(\U1/aes_core/SB3/n1965 ), 
        .B(\U1/aes_core/SB3/n1964 ), .C(\U1/aes_core/SB3/n2043 ), .D(
        \U1/aes_core/SB3/n3266 ), .Y(\U1/aes_core/SB3/n1969 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1156  ( .A(\U1/aes_core/SB3/n3269 ), .B(
        \U1/aes_core/SB3/n3330 ), .Y(\U1/aes_core/SB3/n3313 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1155  ( .AN(\U1/aes_core/SB3/n1967 ), 
        .B(\U1/aes_core/SB3/n1966 ), .C(\U1/aes_core/SB3/n3313 ), .Y(
        \U1/aes_core/SB3/n1968 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1154  ( .A(\U1/aes_core/SB3/n2025 ), .B(
        \U1/aes_core/SB3/n1972 ), .C(\U1/aes_core/SB3/n1971 ), .D(
        \U1/aes_core/SB3/n1970 ), .E(\U1/aes_core/SB3/n1969 ), .F(
        \U1/aes_core/SB3/n1968 ), .Y(\U1/aes_core/SB3/n2001 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1153  ( .A(\U1/aes_core/SB3/n1973 ), .Y(
        \U1/aes_core/SB3/n1975 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1152  ( .A0(\U1/aes_core/SB3/n3322 ), 
        .A1(\U1/aes_core/SB3/n2058 ), .B0(\U1/aes_core/SB3/n2060 ), .B1(
        \U1/aes_core/SB3/n3327 ), .Y(\U1/aes_core/SB3/n1974 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U1151  ( .A0(\U1/aes_core/SB3/n3344 ), 
        .A1(\U1/aes_core/SB3/n3346 ), .B0(\U1/aes_core/SB3/n1975 ), .C0(
        \U1/aes_core/SB3/n1974 ), .Y(\U1/aes_core/SB3/n1986 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1150  ( .A0(\U1/aes_core/SB3/n3324 ), 
        .A1(\U1/aes_core/SB3/n3322 ), .B0(\U1/aes_core/SB3/n2019 ), .Y(
        \U1/aes_core/SB3/n1979 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1149  ( .A0(\U1/aes_core/SB3/n3325 ), 
        .A1(\U1/aes_core/SB3/n3339 ), .B0(\U1/aes_core/SB3/n1976 ), .Y(
        \U1/aes_core/SB3/n1978 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1148  ( .AN(\U1/aes_core/SB3/n1980 ), 
        .B(\U1/aes_core/SB3/n1979 ), .C(\U1/aes_core/SB3/n1978 ), .D(
        \U1/aes_core/SB3/n1977 ), .Y(\U1/aes_core/SB3/n1985 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1147  ( .A0(\U1/aes_core/SB3/n3332 ), 
        .A1(\U1/aes_core/SB3/n3329 ), .B0(\U1/aes_core/SB3/n3333 ), .Y(
        \U1/aes_core/SB3/n1982 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1146  ( .A(\U1/aes_core/SB3/n2017 ), .B(
        \U1/aes_core/SB3/n3302 ), .Y(\U1/aes_core/SB3/n3341 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1145  ( .A0(\U1/aes_core/SB3/n3307 ), 
        .A1(\U1/aes_core/SB3/n3341 ), .B0(\U1/aes_core/SB3/n2054 ), .B1(
        \U1/aes_core/SB3/n3305 ), .Y(\U1/aes_core/SB3/n1981 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U1144  ( .A0(\U1/aes_core/SB3/n1983 ), 
        .A1(\U1/aes_core/SB3/n2039 ), .B0(\U1/aes_core/SB3/n1982 ), .C0(
        \U1/aes_core/SB3/n1981 ), .Y(\U1/aes_core/SB3/n1984 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1143  ( .A(\U1/aes_core/SB3/n2001 ), .B(
        \U1/aes_core/SB3/n1988 ), .C(\U1/aes_core/SB3/n1987 ), .D(
        \U1/aes_core/SB3/n1986 ), .E(\U1/aes_core/SB3/n1985 ), .F(
        \U1/aes_core/SB3/n1984 ), .Y(\U1/aes_core/sb3 [13]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1142  ( .A0(\U1/aes_core/SB3/n3343 ), 
        .A1(\U1/aes_core/SB3/n3296 ), .B0(\U1/aes_core/SB3/n3301 ), .B1(
        \U1/aes_core/SB3/n2070 ), .C0(\U1/aes_core/SB3/n1989 ), .Y(
        \U1/aes_core/SB3/n1998 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1141  ( .A0(\U1/aes_core/SB3/n3275 ), 
        .A1(\U1/aes_core/SB3/n2068 ), .B0(\U1/aes_core/SB3/n3322 ), .Y(
        \U1/aes_core/SB3/n1993 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1140  ( .A0(\U1/aes_core/SB3/n2055 ), 
        .A1(\U1/aes_core/SB3/n3299 ), .B0(\U1/aes_core/SB3/n2060 ), .Y(
        \U1/aes_core/SB3/n1992 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1139  ( .A(\U1/aes_core/SB3/n2010 ), .B(
        \U1/aes_core/SB3/n3346 ), .Y(\U1/aes_core/SB3/n3328 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1138  ( .A0(\U1/aes_core/SB3/n3305 ), 
        .A1(\U1/aes_core/SB3/n3268 ), .B0(\U1/aes_core/SB3/n3328 ), .Y(
        \U1/aes_core/SB3/n1991 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1137  ( .A(\U1/aes_core/SB3/n1993 ), .B(
        \U1/aes_core/SB3/n1992 ), .C(\U1/aes_core/SB3/n1991 ), .D(
        \U1/aes_core/SB3/n1990 ), .Y(\U1/aes_core/SB3/n1997 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1136  ( .A(\U1/aes_core/SB3/n3343 ), .B(
        \U1/aes_core/SB3/n3344 ), .Y(\U1/aes_core/SB3/n2066 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1135  ( .A(\U1/aes_core/SB3/n3332 ), .B(
        \U1/aes_core/SB3/n2066 ), .Y(\U1/aes_core/SB3/n1994 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1134  ( .A0(\U1/aes_core/SB3/n2057 ), 
        .A1(\U1/aes_core/SB3/n1995 ), .B0(\U1/aes_core/SB3/n1994 ), .B1(
        \U1/aes_core/SB3/n2010 ), .C0(\U1/aes_core/SB3/n2008 ), .C1(
        \U1/aes_core/SB3/n2039 ), .Y(\U1/aes_core/SB3/n1996 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1133  ( .A(\U1/aes_core/SB3/n2001 ), .B(
        \U1/aes_core/SB3/n2000 ), .C(\U1/aes_core/SB3/n1999 ), .D(
        \U1/aes_core/SB3/n1998 ), .E(\U1/aes_core/SB3/n1997 ), .F(
        \U1/aes_core/SB3/n1996 ), .Y(\U1/aes_core/sb3 [14]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1132  ( .A0(\U1/aes_core/SB3/n2002 ), 
        .A1(\U1/aes_core/SB3/n3302 ), .B0(\U1/aes_core/SB3/n2070 ), .Y(
        \U1/aes_core/SB3/n2014 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U1131  ( .A(\U1/aes_core/SB3/n2005 ), .B(
        \U1/aes_core/SB3/n2004 ), .C(\U1/aes_core/SB3/n2003 ), .Y(
        \U1/aes_core/SB3/n2013 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U1130  ( .A(\U1/aes_core/SB3/n2054 ), .B(
        \U1/aes_core/SB3/n2058 ), .C(\U1/aes_core/SB3/n3282 ), .Y(
        \U1/aes_core/SB3/n2007 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1129  ( .A0(\U1/aes_core/SB3/n2009 ), 
        .A1(\U1/aes_core/SB3/n2008 ), .B0(\U1/aes_core/SB3/n2007 ), .B1(
        \U1/aes_core/SB3/n2065 ), .C0(\U1/aes_core/SB3/n2006 ), .C1(
        \U1/aes_core/SB3/n3280 ), .Y(\U1/aes_core/SB3/n2012 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U1128  ( .A0(\U1/aes_core/SB3/n3343 ), 
        .A1(\U1/aes_core/SB3/n2039 ), .B0(\U1/aes_core/SB3/n3344 ), .B1(
        \U1/aes_core/SB3/n2010 ), .Y(\U1/aes_core/SB3/n2011 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1127  ( .A(\U1/aes_core/SB3/n2016 ), .B(
        \U1/aes_core/SB3/n2015 ), .C(\U1/aes_core/SB3/n2014 ), .D(
        \U1/aes_core/SB3/n2013 ), .E(\U1/aes_core/SB3/n2012 ), .F(
        \U1/aes_core/SB3/n2011 ), .Y(\U1/aes_core/SB3/n3352 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U1126  ( .A0(\U1/aes_core/SB3/n3278 ), 
        .A1(\U1/aes_core/SB3/n3347 ), .B0(\U1/aes_core/SB3/n2017 ), .Y(
        \U1/aes_core/SB3/n2033 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB3/U1125  ( .A0(\U1/aes_core/SB3/n2019 ), 
        .A1(\U1/aes_core/SB3/n3269 ), .B0(\U1/aes_core/SB3/n2018 ), .B1(
        \U1/aes_core/SB3/n3329 ), .Y(\U1/aes_core/SB3/n2032 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1124  ( .A0(\U1/aes_core/SB3/n3281 ), 
        .A1(\U1/aes_core/SB3/n3344 ), .B0(\U1/aes_core/SB3/n2021 ), .B1(
        \U1/aes_core/SB3/n2020 ), .C0(\U1/aes_core/SB3/n2039 ), .C1(
        \U1/aes_core/SB3/n2065 ), .Y(\U1/aes_core/SB3/n2031 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1123  ( .A(\U1/aes_core/SB3/n2025 ), .B(
        \U1/aes_core/SB3/n2024 ), .C(\U1/aes_core/SB3/n2023 ), .D(
        \U1/aes_core/SB3/n2022 ), .Y(\U1/aes_core/SB3/n2030 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1122  ( .AN(\U1/aes_core/SB3/n2028 ), 
        .B(\U1/aes_core/SB3/n2027 ), .C(\U1/aes_core/SB3/n2026 ), .Y(
        \U1/aes_core/SB3/n2029 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1121  ( .A(\U1/aes_core/SB3/n2034 ), .B(
        \U1/aes_core/SB3/n2033 ), .C(\U1/aes_core/SB3/n2032 ), .D(
        \U1/aes_core/SB3/n2031 ), .E(\U1/aes_core/SB3/n2030 ), .F(
        \U1/aes_core/SB3/n2029 ), .Y(\U1/aes_core/SB3/n3294 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1120  ( .A0(\U1/aes_core/SB3/n3307 ), 
        .A1(\U1/aes_core/SB3/n3327 ), .B0(\U1/aes_core/SB3/n2054 ), .Y(
        \U1/aes_core/SB3/n2038 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1119  ( .A(\U1/aes_core/SB3/n2038 ), .B(
        \U1/aes_core/SB3/n2037 ), .C(\U1/aes_core/SB3/n2036 ), .D(
        \U1/aes_core/SB3/n2035 ), .Y(\U1/aes_core/SB3/n2051 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1118  ( .A0(\U1/aes_core/SB3/n3301 ), 
        .A1(\U1/aes_core/SB3/n2070 ), .B0(\U1/aes_core/SB3/n3279 ), .B1(
        \U1/aes_core/SB3/n3280 ), .C0(\U1/aes_core/SB3/n3309 ), .C1(
        \U1/aes_core/SB3/n2039 ), .Y(\U1/aes_core/SB3/n2050 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1117  ( .A(\U1/aes_core/SB3/n2043 ), .B(
        \U1/aes_core/SB3/n2042 ), .C(\U1/aes_core/SB3/n2041 ), .D(
        \U1/aes_core/SB3/n2040 ), .Y(\U1/aes_core/SB3/n2049 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U1116  ( .A(\U1/aes_core/SB3/n2047 ), .B(
        \U1/aes_core/SB3/n2046 ), .C(\U1/aes_core/SB3/n2045 ), .D(
        \U1/aes_core/SB3/n2044 ), .Y(\U1/aes_core/SB3/n2048 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1115  ( .A(\U1/aes_core/SB3/n2051 ), .B(
        \U1/aes_core/SB3/n2050 ), .C(\U1/aes_core/SB3/n2049 ), .D(
        \U1/aes_core/SB3/n2048 ), .Y(\U1/aes_core/SB3/n2052 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1114  ( .A(\U1/aes_core/SB3/n2052 ), .Y(
        \U1/aes_core/SB3/n3285 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1113  ( .A0(\U1/aes_core/SB3/n2055 ), 
        .A1(\U1/aes_core/SB3/n3330 ), .B0(\U1/aes_core/SB3/n2054 ), .B1(
        \U1/aes_core/SB3/n2053 ), .Y(\U1/aes_core/SB3/n2056 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U1112  ( .A0(\U1/aes_core/SB3/n2057 ), 
        .A1(\U1/aes_core/SB3/n3309 ), .B0(\U1/aes_core/SB3/n3285 ), .C0(
        \U1/aes_core/SB3/n2056 ), .Y(\U1/aes_core/SB3/n2073 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U1111  ( .A1N(\U1/aes_core/SB3/n2059 ), 
        .A0(\U1/aes_core/SB3/n2058 ), .B0(\U1/aes_core/SB3/n3332 ), .Y(
        \U1/aes_core/SB3/n2063 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1110  ( .A0(\U1/aes_core/SB3/n3327 ), 
        .A1(\U1/aes_core/SB3/n3322 ), .B0(\U1/aes_core/SB3/n2060 ), .Y(
        \U1/aes_core/SB3/n2062 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1109  ( .AN(\U1/aes_core/SB3/n2064 ), 
        .B(\U1/aes_core/SB3/n2063 ), .C(\U1/aes_core/SB3/n2062 ), .D(
        \U1/aes_core/SB3/n2061 ), .Y(\U1/aes_core/SB3/n2072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1108  ( .A(\U1/aes_core/SB3/n2065 ), .B(
        \U1/aes_core/SB3/n3343 ), .Y(\U1/aes_core/SB3/n2067 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1107  ( .A0(\U1/aes_core/SB3/n2068 ), 
        .A1(\U1/aes_core/SB3/n2067 ), .B0(\U1/aes_core/SB3/n3282 ), .B1(
        \U1/aes_core/SB3/n2066 ), .Y(\U1/aes_core/SB3/n2069 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1106  ( .A0(\U1/aes_core/SB3/n3281 ), 
        .A1(\U1/aes_core/SB3/n3347 ), .B0(\U1/aes_core/SB3/n2070 ), .B1(
        \U1/aes_core/SB3/n3342 ), .C0(\U1/aes_core/SB3/n2069 ), .Y(
        \U1/aes_core/SB3/n2071 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U1105  ( .A(\U1/aes_core/SB3/n3352 ), .B(
        \U1/aes_core/SB3/n3294 ), .C(\U1/aes_core/SB3/n2074 ), .D(
        \U1/aes_core/SB3/n2073 ), .E(\U1/aes_core/SB3/n2072 ), .F(
        \U1/aes_core/SB3/n2071 ), .Y(\U1/aes_core/sb3 [15]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1104  ( .A(Dout[23]), .B(Dout[22]), .Y(
        \U1/aes_core/SB3/n2093 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1103  ( .A(Dout[21]), .B(Dout[20]), .Y(
        \U1/aes_core/SB3/n2084 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1102  ( .A(\U1/aes_core/SB3/n2093 ), .B(
        \U1/aes_core/SB3/n2084 ), .Y(\U1/aes_core/SB3/n2157 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1101  ( .A(Dout[17]), .Y(
        \U1/aes_core/SB3/n2078 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1100  ( .A(Dout[16]), .Y(
        \U1/aes_core/SB3/n2075 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1099  ( .A(\U1/aes_core/SB3/n2078 ), .B(
        \U1/aes_core/SB3/n2075 ), .Y(\U1/aes_core/SB3/n2085 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1098  ( .A(Dout[19]), .B(Dout[18]), .Y(
        \U1/aes_core/SB3/n2105 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1097  ( .A(\U1/aes_core/SB3/n2085 ), .B(
        \U1/aes_core/SB3/n2105 ), .Y(\U1/aes_core/SB3/n2464 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1096  ( .A(\U1/aes_core/SB3/n2157 ), .B(
        \U1/aes_core/SB3/n2464 ), .Y(\U1/aes_core/SB3/n2246 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U1095  ( .A(Dout[18]), .B(Dout[19]), .Y(
        \U1/aes_core/SB3/n2088 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1094  ( .A(\U1/aes_core/SB3/n2088 ), .B(
        \U1/aes_core/SB3/n2085 ), .Y(\U1/aes_core/SB3/n2402 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1093  ( .A(Dout[23]), .Y(
        \U1/aes_core/SB3/n2081 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1092  ( .A(\U1/aes_core/SB3/n2081 ), .B(
        Dout[22]), .Y(\U1/aes_core/SB3/n2111 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1091  ( .A(\U1/aes_core/SB3/n2111 ), .B(
        \U1/aes_core/SB3/n2084 ), .Y(\U1/aes_core/SB3/n2156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1090  ( .A(\U1/aes_core/SB3/n2402 ), .B(
        \U1/aes_core/SB3/n2156 ), .Y(\U1/aes_core/SB3/n2368 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1089  ( .A(Dout[19]), .Y(
        \U1/aes_core/SB3/n2076 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U1088  ( .A(Dout[18]), .B(
        \U1/aes_core/SB3/n2076 ), .Y(\U1/aes_core/SB3/n2086 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1087  ( .A(\U1/aes_core/SB3/n2085 ), .B(
        \U1/aes_core/SB3/n2086 ), .Y(\U1/aes_core/SB3/n2308 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1086  ( .A(\U1/aes_core/SB3/n2308 ), .Y(
        \U1/aes_core/SB3/n2498 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1085  ( .A(Dout[20]), .Y(
        \U1/aes_core/SB3/n2077 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1084  ( .A(\U1/aes_core/SB3/n2077 ), .B(
        Dout[21]), .Y(\U1/aes_core/SB3/n2092 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1083  ( .A(Dout[22]), .Y(
        \U1/aes_core/SB3/n2080 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1082  ( .A(\U1/aes_core/SB3/n2080 ), .B(
        Dout[23]), .Y(\U1/aes_core/SB3/n2102 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1081  ( .A(\U1/aes_core/SB3/n2092 ), .B(
        \U1/aes_core/SB3/n2102 ), .Y(\U1/aes_core/SB3/n2354 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1080  ( .A(\U1/aes_core/SB3/n2354 ), .Y(
        \U1/aes_core/SB3/n2452 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1079  ( .A(\U1/aes_core/SB3/n2498 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2286 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1078  ( .A(\U1/aes_core/SB3/n2157 ), .Y(
        \U1/aes_core/SB3/n2467 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1077  ( .A(Dout[17]), .B(Dout[16]), .Y(
        \U1/aes_core/SB3/n2089 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1076  ( .A(\U1/aes_core/SB3/n2089 ), .B(
        \U1/aes_core/SB3/n2105 ), .Y(\U1/aes_core/SB3/n2420 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1075  ( .A(\U1/aes_core/SB3/n2420 ), .Y(
        \U1/aes_core/SB3/n2508 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1074  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2508 ), .Y(\U1/aes_core/SB3/n2425 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1073  ( .A(\U1/aes_core/SB3/n2075 ), .B(
        Dout[17]), .Y(\U1/aes_core/SB3/n2104 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1072  ( .A(\U1/aes_core/SB3/n2086 ), .B(
        \U1/aes_core/SB3/n2104 ), .Y(\U1/aes_core/SB3/n2295 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1071  ( .A(\U1/aes_core/SB3/n2295 ), .Y(
        \U1/aes_core/SB3/n2409 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1070  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2264 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U1069  ( .A(\U1/aes_core/SB3/n2286 ), .B(
        \U1/aes_core/SB3/n2425 ), .C(\U1/aes_core/SB3/n2264 ), .Y(
        \U1/aes_core/SB3/n2124 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1068  ( .A(\U1/aes_core/SB3/n2084 ), .B(
        \U1/aes_core/SB3/n2102 ), .Y(\U1/aes_core/SB3/n2353 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1067  ( .A(\U1/aes_core/SB3/n2076 ), .B(
        Dout[18]), .Y(\U1/aes_core/SB3/n2095 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1066  ( .A(\U1/aes_core/SB3/n2095 ), .B(
        \U1/aes_core/SB3/n2104 ), .Y(\U1/aes_core/SB3/n2351 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1065  ( .A(\U1/aes_core/SB3/n2353 ), .B(
        \U1/aes_core/SB3/n2351 ), .Y(\U1/aes_core/SB3/n2241 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1064  ( .A(\U1/aes_core/SB3/n2156 ), .Y(
        \U1/aes_core/SB3/n2469 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1063  ( .A(Dout[21]), .Y(
        \U1/aes_core/SB3/n2079 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1062  ( .A(\U1/aes_core/SB3/n2077 ), .B(
        \U1/aes_core/SB3/n2079 ), .Y(\U1/aes_core/SB3/n2103 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1061  ( .A(\U1/aes_core/SB3/n2093 ), .B(
        \U1/aes_core/SB3/n2103 ), .Y(\U1/aes_core/SB3/n2512 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1060  ( .A(\U1/aes_core/SB3/n2512 ), .Y(
        \U1/aes_core/SB3/n2443 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1059  ( .A(\U1/aes_core/SB3/n2078 ), .B(
        Dout[16]), .Y(\U1/aes_core/SB3/n2094 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1058  ( .A(\U1/aes_core/SB3/n2094 ), .B(
        \U1/aes_core/SB3/n2105 ), .Y(\U1/aes_core/SB3/n2477 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1057  ( .A(\U1/aes_core/SB3/n2477 ), .Y(
        \U1/aes_core/SB3/n2300 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1056  ( .A0(\U1/aes_core/SB3/n2469 ), 
        .A1(\U1/aes_core/SB3/n2443 ), .B0(\U1/aes_core/SB3/n2300 ), .Y(
        \U1/aes_core/SB3/n2083 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1055  ( .A(\U1/aes_core/SB3/n2089 ), .B(
        \U1/aes_core/SB3/n2086 ), .Y(\U1/aes_core/SB3/n2465 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1054  ( .A(\U1/aes_core/SB3/n2465 ), .Y(
        \U1/aes_core/SB3/n2451 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1053  ( .A(\U1/aes_core/SB3/n2079 ), .B(
        Dout[20]), .Y(\U1/aes_core/SB3/n2110 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1052  ( .A(\U1/aes_core/SB3/n2102 ), .B(
        \U1/aes_core/SB3/n2110 ), .Y(\U1/aes_core/SB3/n2505 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1051  ( .A(\U1/aes_core/SB3/n2353 ), .B(
        \U1/aes_core/SB3/n2505 ), .Y(\U1/aes_core/SB3/n2219 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1050  ( .A(\U1/aes_core/SB3/n2081 ), .B(
        \U1/aes_core/SB3/n2080 ), .Y(\U1/aes_core/SB3/n2101 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1049  ( .A(\U1/aes_core/SB3/n2092 ), .B(
        \U1/aes_core/SB3/n2101 ), .Y(\U1/aes_core/SB3/n2480 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1048  ( .A(\U1/aes_core/SB3/n2480 ), .Y(
        \U1/aes_core/SB3/n2200 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1047  ( .A0(\U1/aes_core/SB3/n2451 ), 
        .A1(\U1/aes_core/SB3/n2219 ), .B0(\U1/aes_core/SB3/n2200 ), .B1(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2082 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U1046  ( .AN(\U1/aes_core/SB3/n2241 ), 
        .B(\U1/aes_core/SB3/n2083 ), .C(\U1/aes_core/SB3/n2082 ), .Y(
        \U1/aes_core/SB3/n2123 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1045  ( .A(\U1/aes_core/SB3/n2084 ), .B(
        \U1/aes_core/SB3/n2101 ), .Y(\U1/aes_core/SB3/n2370 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1044  ( .A(\U1/aes_core/SB3/n2088 ), .B(
        \U1/aes_core/SB3/n2089 ), .Y(\U1/aes_core/SB3/n2515 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1043  ( .A(\U1/aes_core/SB3/n2111 ), .B(
        \U1/aes_core/SB3/n2092 ), .Y(\U1/aes_core/SB3/n2421 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1042  ( .A(\U1/aes_core/SB3/n2088 ), .B(
        \U1/aes_core/SB3/n2094 ), .Y(\U1/aes_core/SB3/n2418 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1041  ( .A(\U1/aes_core/SB3/n2085 ), .B(
        \U1/aes_core/SB3/n2095 ), .Y(\U1/aes_core/SB3/n2423 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1040  ( .A(\U1/aes_core/SB3/n2423 ), .Y(
        \U1/aes_core/SB3/n2403 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1039  ( .A(\U1/aes_core/SB3/n2505 ), .Y(
        \U1/aes_core/SB3/n2214 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1038  ( .A(\U1/aes_core/SB3/n2086 ), .B(
        \U1/aes_core/SB3/n2094 ), .Y(\U1/aes_core/SB3/n2441 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1037  ( .A(\U1/aes_core/SB3/n2441 ), .Y(
        \U1/aes_core/SB3/n2466 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U1036  ( .A0(\U1/aes_core/SB3/n2403 ), 
        .A1(\U1/aes_core/SB3/n2467 ), .B0(\U1/aes_core/SB3/n2214 ), .B1(
        \U1/aes_core/SB3/n2466 ), .Y(\U1/aes_core/SB3/n2087 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U1035  ( .A0(\U1/aes_core/SB3/n2370 ), 
        .A1(\U1/aes_core/SB3/n2515 ), .B0(\U1/aes_core/SB3/n2421 ), .B1(
        \U1/aes_core/SB3/n2418 ), .C0(\U1/aes_core/SB3/n2087 ), .Y(
        \U1/aes_core/SB3/n2122 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1034  ( .A(\U1/aes_core/SB3/n2423 ), .B(
        \U1/aes_core/SB3/n2370 ), .Y(\U1/aes_core/SB3/n2207 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1033  ( .A(\U1/aes_core/SB3/n2418 ), .B(
        \U1/aes_core/SB3/n2353 ), .Y(\U1/aes_core/SB3/n2217 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1032  ( .A(\U1/aes_core/SB3/n2217 ), .Y(
        \U1/aes_core/SB3/n2091 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1031  ( .A(\U1/aes_core/SB3/n2088 ), .B(
        \U1/aes_core/SB3/n2104 ), .Y(\U1/aes_core/SB3/n2493 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1030  ( .A(\U1/aes_core/SB3/n2493 ), .Y(
        \U1/aes_core/SB3/n2442 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1029  ( .A(\U1/aes_core/SB3/n2089 ), .B(
        \U1/aes_core/SB3/n2095 ), .Y(\U1/aes_core/SB3/n2478 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1028  ( .A(\U1/aes_core/SB3/n2478 ), .Y(
        \U1/aes_core/SB3/n2489 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U1027  ( .A0(\U1/aes_core/SB3/n2442 ), 
        .A1(\U1/aes_core/SB3/n2489 ), .B0(\U1/aes_core/SB3/n2443 ), .Y(
        \U1/aes_core/SB3/n2090 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1026  ( .A(\U1/aes_core/SB3/n2093 ), .B(
        \U1/aes_core/SB3/n2110 ), .Y(\U1/aes_core/SB3/n2494 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1025  ( .A(\U1/aes_core/SB3/n2494 ), .Y(
        \U1/aes_core/SB3/n2444 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1024  ( .A(\U1/aes_core/SB3/n2444 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2234 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1023  ( .AN(\U1/aes_core/SB3/n2207 ), 
        .B(\U1/aes_core/SB3/n2091 ), .C(\U1/aes_core/SB3/n2090 ), .D(
        \U1/aes_core/SB3/n2234 ), .Y(\U1/aes_core/SB3/n2100 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1022  ( .A(\U1/aes_core/SB3/n2103 ), .B(
        \U1/aes_core/SB3/n2101 ), .Y(\U1/aes_core/SB3/n2514 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1021  ( .A(\U1/aes_core/SB3/n2093 ), .B(
        \U1/aes_core/SB3/n2092 ), .Y(\U1/aes_core/SB3/n2506 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U1020  ( .A0(\U1/aes_core/SB3/n2156 ), 
        .A1(\U1/aes_core/SB3/n2308 ), .B0(\U1/aes_core/SB3/n2514 ), .B1(
        \U1/aes_core/SB3/n2423 ), .C0(\U1/aes_core/SB3/n2506 ), .C1(
        \U1/aes_core/SB3/n2441 ), .Y(\U1/aes_core/SB3/n2099 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1019  ( .A(\U1/aes_core/SB3/n2465 ), .B(
        \U1/aes_core/SB3/n2156 ), .Y(\U1/aes_core/SB3/n2292 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1018  ( .A(\U1/aes_core/SB3/n2214 ), .B(
        \U1/aes_core/SB3/n2403 ), .Y(\U1/aes_core/SB3/n2245 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1017  ( .A(\U1/aes_core/SB3/n2466 ), .B(
        \U1/aes_core/SB3/n2467 ), .Y(\U1/aes_core/SB3/n2265 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1016  ( .A(\U1/aes_core/SB3/n2421 ), .Y(
        \U1/aes_core/SB3/n2495 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1015  ( .A(\U1/aes_core/SB3/n2495 ), .B(
        \U1/aes_core/SB3/n2300 ), .Y(\U1/aes_core/SB3/n2303 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1014  ( .AN(\U1/aes_core/SB3/n2292 ), 
        .B(\U1/aes_core/SB3/n2245 ), .C(\U1/aes_core/SB3/n2265 ), .D(
        \U1/aes_core/SB3/n2303 ), .Y(\U1/aes_core/SB3/n2098 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1013  ( .A(\U1/aes_core/SB3/n2111 ), .B(
        \U1/aes_core/SB3/n2103 ), .Y(\U1/aes_core/SB3/n2215 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1012  ( .A(\U1/aes_core/SB3/n2215 ), .B(
        \U1/aes_core/SB3/n2477 ), .Y(\U1/aes_core/SB3/n2394 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1011  ( .A(\U1/aes_core/SB3/n2095 ), .B(
        \U1/aes_core/SB3/n2094 ), .Y(\U1/aes_core/SB3/n2513 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1010  ( .A(\U1/aes_core/SB3/n2480 ), .B(
        \U1/aes_core/SB3/n2513 ), .Y(\U1/aes_core/SB3/n2359 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1009  ( .A(\U1/aes_core/SB3/n2359 ), .Y(
        \U1/aes_core/SB3/n2096 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1008  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2300 ), .Y(\U1/aes_core/SB3/n2378 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1007  ( .A(\U1/aes_core/SB3/n2513 ), .Y(
        \U1/aes_core/SB3/n2496 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1006  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2496 ), .Y(\U1/aes_core/SB3/n2429 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U1005  ( .AN(\U1/aes_core/SB3/n2394 ), 
        .B(\U1/aes_core/SB3/n2096 ), .C(\U1/aes_core/SB3/n2378 ), .D(
        \U1/aes_core/SB3/n2429 ), .Y(\U1/aes_core/SB3/n2097 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U1004  ( .A(\U1/aes_core/SB3/n2100 ), .B(
        \U1/aes_core/SB3/n2099 ), .C(\U1/aes_core/SB3/n2098 ), .D(
        \U1/aes_core/SB3/n2097 ), .Y(\U1/aes_core/SB3/n2196 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1003  ( .A(\U1/aes_core/SB3/n2420 ), .B(
        \U1/aes_core/SB3/n2215 ), .Y(\U1/aes_core/SB3/n2428 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U1002  ( .A(\U1/aes_core/SB3/n2110 ), .B(
        \U1/aes_core/SB3/n2101 ), .Y(\U1/aes_core/SB3/n2311 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U1001  ( .A(\U1/aes_core/SB3/n2402 ), .B(
        \U1/aes_core/SB3/n2311 ), .Y(\U1/aes_core/SB3/n2282 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U1000  ( .A(\U1/aes_core/SB3/n2514 ), .Y(
        \U1/aes_core/SB3/n2470 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U999  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2451 ), .Y(\U1/aes_core/SB3/n2231 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U998  ( .A0(\U1/aes_core/SB3/n2311 ), 
        .A1(\U1/aes_core/SB3/n2513 ), .B0(\U1/aes_core/SB3/n2231 ), .Y(
        \U1/aes_core/SB3/n2109 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U997  ( .A(\U1/aes_core/SB3/n2351 ), .Y(
        \U1/aes_core/SB3/n2446 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U996  ( .A(\U1/aes_core/SB3/n2446 ), .B(
        \U1/aes_core/SB3/n2469 ), .Y(\U1/aes_core/SB3/n2447 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U995  ( .A(\U1/aes_core/SB3/n2469 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2406 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U994  ( .A(\U1/aes_core/SB3/n2103 ), .B(
        \U1/aes_core/SB3/n2102 ), .Y(\U1/aes_core/SB3/n2476 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U993  ( .A(\U1/aes_core/SB3/n2476 ), .Y(
        \U1/aes_core/SB3/n2226 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U992  ( .A(\U1/aes_core/SB3/n2442 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2250 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U991  ( .A(\U1/aes_core/SB3/n2464 ), .Y(
        \U1/aes_core/SB3/n2445 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U990  ( .A(\U1/aes_core/SB3/n2445 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2314 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U989  ( .A(\U1/aes_core/SB3/n2447 ), .B(
        \U1/aes_core/SB3/n2406 ), .C(\U1/aes_core/SB3/n2250 ), .D(
        \U1/aes_core/SB3/n2314 ), .Y(\U1/aes_core/SB3/n2108 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U988  ( .A(\U1/aes_core/SB3/n2466 ), .B(
        \U1/aes_core/SB3/n2444 ), .Y(\U1/aes_core/SB3/n2373 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U987  ( .A(\U1/aes_core/SB3/n2508 ), .B(
        \U1/aes_core/SB3/n2444 ), .Y(\U1/aes_core/SB3/n2364 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U986  ( .A(\U1/aes_core/SB3/n2506 ), .Y(
        \U1/aes_core/SB3/n2499 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U985  ( .A(\U1/aes_core/SB3/n2403 ), .B(
        \U1/aes_core/SB3/n2499 ), .Y(\U1/aes_core/SB3/n2211 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U984  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2442 ), .Y(\U1/aes_core/SB3/n2347 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U983  ( .A(\U1/aes_core/SB3/n2373 ), .B(
        \U1/aes_core/SB3/n2364 ), .C(\U1/aes_core/SB3/n2211 ), .D(
        \U1/aes_core/SB3/n2347 ), .Y(\U1/aes_core/SB3/n2107 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U982  ( .A(\U1/aes_core/SB3/n2418 ), .Y(
        \U1/aes_core/SB3/n2387 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U981  ( .A(\U1/aes_core/SB3/n2214 ), .B(
        \U1/aes_core/SB3/n2387 ), .Y(\U1/aes_core/SB3/n2198 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U980  ( .A(\U1/aes_core/SB3/n2105 ), .B(
        \U1/aes_core/SB3/n2104 ), .Y(\U1/aes_core/SB3/n2453 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U979  ( .A(\U1/aes_core/SB3/n2453 ), .Y(
        \U1/aes_core/SB3/n2487 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U978  ( .A(\U1/aes_core/SB3/n2214 ), .B(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2262 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U977  ( .A(\U1/aes_core/SB3/n2402 ), .Y(
        \U1/aes_core/SB3/n2510 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U976  ( .A(\U1/aes_core/SB3/n2510 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2297 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U975  ( .A(\U1/aes_core/SB3/n2443 ), .B(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2471 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U974  ( .A(\U1/aes_core/SB3/n2198 ), .B(
        \U1/aes_core/SB3/n2262 ), .C(\U1/aes_core/SB3/n2297 ), .D(
        \U1/aes_core/SB3/n2471 ), .Y(\U1/aes_core/SB3/n2106 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U973  ( .A(\U1/aes_core/SB3/n2428 ), .B(
        \U1/aes_core/SB3/n2282 ), .C(\U1/aes_core/SB3/n2109 ), .D(
        \U1/aes_core/SB3/n2108 ), .E(\U1/aes_core/SB3/n2107 ), .F(
        \U1/aes_core/SB3/n2106 ), .Y(\U1/aes_core/SB3/n2185 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U972  ( .A(\U1/aes_core/SB3/n2185 ), .Y(
        \U1/aes_core/SB3/n2120 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U971  ( .A(\U1/aes_core/SB3/n2478 ), .B(
        \U1/aes_core/SB3/n2311 ), .Y(\U1/aes_core/SB3/n2208 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U970  ( .A(\U1/aes_core/SB3/n2111 ), .B(
        \U1/aes_core/SB3/n2110 ), .Y(\U1/aes_core/SB3/n2475 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U969  ( .A(\U1/aes_core/SB3/n2475 ), .B(
        \U1/aes_core/SB3/n2351 ), .Y(\U1/aes_core/SB3/n2360 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U968  ( .A(\U1/aes_core/SB3/n2360 ), .Y(
        \U1/aes_core/SB3/n2113 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U967  ( .A(\U1/aes_core/SB3/n2353 ), .Y(
        \U1/aes_core/SB3/n2500 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U966  ( .A0(\U1/aes_core/SB3/n2226 ), 
        .A1(\U1/aes_core/SB3/n2500 ), .B0(\U1/aes_core/SB3/n2487 ), .Y(
        \U1/aes_core/SB3/n2112 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U965  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2387 ), .Y(\U1/aes_core/SB3/n2233 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U964  ( .AN(\U1/aes_core/SB3/n2208 ), 
        .B(\U1/aes_core/SB3/n2113 ), .C(\U1/aes_core/SB3/n2112 ), .D(
        \U1/aes_core/SB3/n2233 ), .Y(\U1/aes_core/SB3/n2117 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U963  ( .A0(\U1/aes_core/SB3/n2464 ), 
        .A1(\U1/aes_core/SB3/n2512 ), .B0(\U1/aes_core/SB3/n2370 ), .B1(
        \U1/aes_core/SB3/n2418 ), .C0(\U1/aes_core/SB3/n2477 ), .C1(
        \U1/aes_core/SB3/n2494 ), .Y(\U1/aes_core/SB3/n2116 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U962  ( .A(\U1/aes_core/SB3/n2512 ), .B(
        \U1/aes_core/SB3/n2515 ), .Y(\U1/aes_core/SB3/n2273 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U961  ( .A(\U1/aes_core/SB3/n2500 ), .B(
        \U1/aes_core/SB3/n2442 ), .Y(\U1/aes_core/SB3/n2431 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U960  ( .A(\U1/aes_core/SB3/n2403 ), .B(
        \U1/aes_core/SB3/n2500 ), .Y(\U1/aes_core/SB3/n2365 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U959  ( .A(\U1/aes_core/SB3/n2387 ), .B(
        \U1/aes_core/SB3/n2467 ), .Y(\U1/aes_core/SB3/n2212 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U958  ( .AN(\U1/aes_core/SB3/n2273 ), 
        .B(\U1/aes_core/SB3/n2431 ), .C(\U1/aes_core/SB3/n2365 ), .D(
        \U1/aes_core/SB3/n2212 ), .Y(\U1/aes_core/SB3/n2115 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U957  ( .A(\U1/aes_core/SB3/n2510 ), .B(
        \U1/aes_core/SB3/n2495 ), .Y(\U1/aes_core/SB3/n2285 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U956  ( .A(\U1/aes_core/SB3/n2387 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2377 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U955  ( .A(\U1/aes_core/SB3/n2214 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2253 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U954  ( .A(\U1/aes_core/SB3/n2446 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2298 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U953  ( .A(\U1/aes_core/SB3/n2285 ), .B(
        \U1/aes_core/SB3/n2377 ), .C(\U1/aes_core/SB3/n2253 ), .D(
        \U1/aes_core/SB3/n2298 ), .Y(\U1/aes_core/SB3/n2114 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U952  ( .A(\U1/aes_core/SB3/n2117 ), .B(
        \U1/aes_core/SB3/n2116 ), .C(\U1/aes_core/SB3/n2115 ), .D(
        \U1/aes_core/SB3/n2114 ), .Y(\U1/aes_core/SB3/n2118 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U951  ( .A(\U1/aes_core/SB3/n2118 ), .Y(
        \U1/aes_core/SB3/n2492 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U950  ( .A(\U1/aes_core/SB3/n2508 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2119 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U949  ( .AN(\U1/aes_core/SB3/n2196 ), 
        .B(\U1/aes_core/SB3/n2120 ), .C(\U1/aes_core/SB3/n2492 ), .D(
        \U1/aes_core/SB3/n2119 ), .Y(\U1/aes_core/SB3/n2121 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U948  ( .A(\U1/aes_core/SB3/n2246 ), .B(
        \U1/aes_core/SB3/n2368 ), .C(\U1/aes_core/SB3/n2124 ), .D(
        \U1/aes_core/SB3/n2123 ), .E(\U1/aes_core/SB3/n2122 ), .F(
        \U1/aes_core/SB3/n2121 ), .Y(\U1/aes_core/SB3/n2175 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U947  ( .A(\U1/aes_core/SB3/n2493 ), .B(
        \U1/aes_core/SB3/n2156 ), .Y(\U1/aes_core/SB3/n2291 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U946  ( .A(\U1/aes_core/SB3/n2443 ), .B(
        \U1/aes_core/SB3/n2510 ), .Y(\U1/aes_core/SB3/n2367 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U945  ( .A(\U1/aes_core/SB3/n2499 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2244 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U944  ( .A(\U1/aes_core/SB3/n2215 ), .Y(
        \U1/aes_core/SB3/n2488 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U943  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2267 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U942  ( .AN(\U1/aes_core/SB3/n2291 ), 
        .B(\U1/aes_core/SB3/n2367 ), .C(\U1/aes_core/SB3/n2244 ), .D(
        \U1/aes_core/SB3/n2267 ), .Y(\U1/aes_core/SB3/n2131 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U941  ( .A(\U1/aes_core/SB3/n2480 ), .B(
        \U1/aes_core/SB3/n2351 ), .Y(\U1/aes_core/SB3/n2393 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U940  ( .A(\U1/aes_core/SB3/n2403 ), .B(
        \U1/aes_core/SB3/n2469 ), .Y(\U1/aes_core/SB3/n2224 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U939  ( .A0(\U1/aes_core/SB3/n2489 ), 
        .A1(\U1/aes_core/SB3/n2409 ), .B0(\U1/aes_core/SB3/n2214 ), .Y(
        \U1/aes_core/SB3/n2125 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U938  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2316 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U937  ( .AN(\U1/aes_core/SB3/n2393 ), 
        .B(\U1/aes_core/SB3/n2224 ), .C(\U1/aes_core/SB3/n2125 ), .D(
        \U1/aes_core/SB3/n2316 ), .Y(\U1/aes_core/SB3/n2126 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U936  ( .A(\U1/aes_core/SB3/n2126 ), .Y(
        \U1/aes_core/SB3/n2130 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U935  ( .A(\U1/aes_core/SB3/n2370 ), .Y(
        \U1/aes_core/SB3/n2490 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U934  ( .A(\U1/aes_core/SB3/n2515 ), .Y(
        \U1/aes_core/SB3/n2410 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U933  ( .A0(\U1/aes_core/SB3/n2510 ), 
        .A1(\U1/aes_core/SB3/n2444 ), .B0(\U1/aes_core/SB3/n2490 ), .B1(
        \U1/aes_core/SB3/n2300 ), .C0(\U1/aes_core/SB3/n2410 ), .C1(
        \U1/aes_core/SB3/n2488 ), .Y(\U1/aes_core/SB3/n2129 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U932  ( .A0(\U1/aes_core/SB3/n2311 ), 
        .A1(\U1/aes_core/SB3/n2493 ), .B0(\U1/aes_core/SB3/n2513 ), .B1(
        \U1/aes_core/SB3/n2514 ), .Y(\U1/aes_core/SB3/n2127 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U931  ( .A0(\U1/aes_core/SB3/n2387 ), 
        .A1(\U1/aes_core/SB3/n2200 ), .B0(\U1/aes_core/SB3/n2443 ), .B1(
        \U1/aes_core/SB3/n2466 ), .C0(\U1/aes_core/SB3/n2127 ), .Y(
        \U1/aes_core/SB3/n2128 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U930  ( .AN(\U1/aes_core/SB3/n2131 ), 
        .B(\U1/aes_core/SB3/n2130 ), .C(\U1/aes_core/SB3/n2129 ), .D(
        \U1/aes_core/SB3/n2128 ), .Y(\U1/aes_core/SB3/n2194 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U929  ( .A(\U1/aes_core/SB3/n2514 ), .B(
        \U1/aes_core/SB3/n2351 ), .Y(\U1/aes_core/SB3/n2209 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U928  ( .A0(\U1/aes_core/SB3/n2421 ), 
        .A1(\U1/aes_core/SB3/n2514 ), .B0(\U1/aes_core/SB3/n2453 ), .Y(
        \U1/aes_core/SB3/n2136 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U927  ( .A(\U1/aes_core/SB3/n2453 ), .B(
        \U1/aes_core/SB3/n2441 ), .Y(\U1/aes_core/SB3/n2293 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB3/U926  ( .A0(\U1/aes_core/SB3/n2442 ), .A1(
        \U1/aes_core/SB3/n2200 ), .B0(\U1/aes_core/SB3/n2293 ), .B1(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2135 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U925  ( .A0(\U1/aes_core/SB3/n2475 ), 
        .A1(\U1/aes_core/SB3/n2515 ), .B0(\U1/aes_core/SB3/n2215 ), .B1(
        \U1/aes_core/SB3/n2308 ), .C0(\U1/aes_core/SB3/n2477 ), .C1(
        \U1/aes_core/SB3/n2506 ), .Y(\U1/aes_core/SB3/n2134 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U924  ( .A(\U1/aes_core/SB3/n2311 ), .Y(
        \U1/aes_core/SB3/n2404 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U923  ( .A(\U1/aes_core/SB3/n2508 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2430 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U922  ( .A(\U1/aes_core/SB3/n2403 ), .B(
        \U1/aes_core/SB3/n2200 ), .Y(\U1/aes_core/SB3/n2232 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U921  ( .A(\U1/aes_core/SB3/n2214 ), .B(
        \U1/aes_core/SB3/n2446 ), .Y(\U1/aes_core/SB3/n2252 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U920  ( .A(\U1/aes_core/SB3/n2403 ), .B(
        \U1/aes_core/SB3/n2444 ), .Y(\U1/aes_core/SB3/n2376 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U919  ( .A(\U1/aes_core/SB3/n2430 ), .B(
        \U1/aes_core/SB3/n2232 ), .C(\U1/aes_core/SB3/n2252 ), .D(
        \U1/aes_core/SB3/n2376 ), .Y(\U1/aes_core/SB3/n2133 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U918  ( .A(\U1/aes_core/SB3/n2423 ), .B(
        \U1/aes_core/SB3/n2311 ), .Y(\U1/aes_core/SB3/n2274 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U917  ( .A(\U1/aes_core/SB3/n2409 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2284 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U916  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2300 ), .Y(\U1/aes_core/SB3/n2315 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U915  ( .AN(\U1/aes_core/SB3/n2274 ), 
        .B(\U1/aes_core/SB3/n2284 ), .C(\U1/aes_core/SB3/n2315 ), .Y(
        \U1/aes_core/SB3/n2132 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U914  ( .A(\U1/aes_core/SB3/n2209 ), .B(
        \U1/aes_core/SB3/n2136 ), .C(\U1/aes_core/SB3/n2135 ), .D(
        \U1/aes_core/SB3/n2134 ), .E(\U1/aes_core/SB3/n2133 ), .F(
        \U1/aes_core/SB3/n2132 ), .Y(\U1/aes_core/SB3/n2521 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U913  ( .A0(\U1/aes_core/SB3/n2214 ), 
        .A1(\U1/aes_core/SB3/n2467 ), .B0(\U1/aes_core/SB3/n2498 ), .Y(
        \U1/aes_core/SB3/n2137 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U912  ( .A(\U1/aes_core/SB3/n2200 ), .B(
        \U1/aes_core/SB3/n2300 ), .Y(\U1/aes_core/SB3/n2362 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U911  ( .A(\U1/aes_core/SB3/n2442 ), .B(
        \U1/aes_core/SB3/n2490 ), .Y(\U1/aes_core/SB3/n2229 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U910  ( .A(\U1/aes_core/SB3/n2490 ), .B(
        \U1/aes_core/SB3/n2446 ), .Y(\U1/aes_core/SB3/n2280 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U909  ( .A(\U1/aes_core/SB3/n2137 ), .B(
        \U1/aes_core/SB3/n2362 ), .C(\U1/aes_core/SB3/n2229 ), .D(
        \U1/aes_core/SB3/n2280 ), .Y(\U1/aes_core/SB3/n2141 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U908  ( .A0(\U1/aes_core/SB3/n2493 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2215 ), .B1(
        \U1/aes_core/SB3/n2465 ), .C0(\U1/aes_core/SB3/n2494 ), .C1(
        \U1/aes_core/SB3/n2351 ), .Y(\U1/aes_core/SB3/n2140 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U907  ( .A(\U1/aes_core/SB3/n2445 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2261 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U906  ( .A(\U1/aes_core/SB3/n2444 ), .B(
        \U1/aes_core/SB3/n2496 ), .Y(\U1/aes_core/SB3/n2426 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U905  ( .A(\U1/aes_core/SB3/n2444 ), .B(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2248 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U904  ( .A(\U1/aes_core/SB3/n2499 ), .B(
        \U1/aes_core/SB3/n2489 ), .Y(\U1/aes_core/SB3/n2210 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U903  ( .A(\U1/aes_core/SB3/n2261 ), .B(
        \U1/aes_core/SB3/n2426 ), .C(\U1/aes_core/SB3/n2248 ), .D(
        \U1/aes_core/SB3/n2210 ), .Y(\U1/aes_core/SB3/n2139 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U902  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2348 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U901  ( .A(\U1/aes_core/SB3/n2508 ), .B(
        \U1/aes_core/SB3/n2469 ), .Y(\U1/aes_core/SB3/n2296 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U900  ( .A(\U1/aes_core/SB3/n2498 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2372 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U899  ( .A(\U1/aes_core/SB3/n2226 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2197 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U898  ( .A(\U1/aes_core/SB3/n2348 ), .B(
        \U1/aes_core/SB3/n2296 ), .C(\U1/aes_core/SB3/n2372 ), .D(
        \U1/aes_core/SB3/n2197 ), .Y(\U1/aes_core/SB3/n2138 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U897  ( .A(\U1/aes_core/SB3/n2141 ), .B(
        \U1/aes_core/SB3/n2140 ), .C(\U1/aes_core/SB3/n2139 ), .D(
        \U1/aes_core/SB3/n2138 ), .Y(\U1/aes_core/SB3/n2183 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U896  ( .A(\U1/aes_core/SB3/n2175 ), .B(
        \U1/aes_core/SB3/n2194 ), .C(\U1/aes_core/SB3/n2521 ), .D(
        \U1/aes_core/SB3/n2183 ), .Y(\U1/aes_core/SB3/n2150 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U895  ( .A(\U1/aes_core/SB3/n2475 ), .Y(
        \U1/aes_core/SB3/n2399 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U894  ( .A0(\U1/aes_core/SB3/n2351 ), 
        .A1(\U1/aes_core/SB3/n2157 ), .B0(\U1/aes_core/SB3/n2295 ), .B1(
        \U1/aes_core/SB3/n2506 ), .Y(\U1/aes_core/SB3/n2142 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U893  ( .A0(\U1/aes_core/SB3/n2399 ), 
        .A1(\U1/aes_core/SB3/n2451 ), .B0(\U1/aes_core/SB3/n2500 ), .B1(
        \U1/aes_core/SB3/n2508 ), .C0(\U1/aes_core/SB3/n2142 ), .Y(
        \U1/aes_core/SB3/n2149 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U892  ( .A(\U1/aes_core/SB3/n2420 ), .B(
        \U1/aes_core/SB3/n2423 ), .Y(\U1/aes_core/SB3/n2419 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U891  ( .A0(\U1/aes_core/SB3/n2354 ), 
        .A1(\U1/aes_core/SB3/n2423 ), .B0(\U1/aes_core/SB3/n2311 ), .B1(
        \U1/aes_core/SB3/n2464 ), .Y(\U1/aes_core/SB3/n2143 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U890  ( .A0(\U1/aes_core/SB3/n2226 ), 
        .A1(\U1/aes_core/SB3/n2419 ), .B0(\U1/aes_core/SB3/n2470 ), .B1(
        \U1/aes_core/SB3/n2489 ), .C0(\U1/aes_core/SB3/n2143 ), .Y(
        \U1/aes_core/SB3/n2148 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U889  ( .A(\U1/aes_core/SB3/n2494 ), .B(
        \U1/aes_core/SB3/n2353 ), .Y(\U1/aes_core/SB3/n2146 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U888  ( .A(\U1/aes_core/SB3/n2444 ), .B(
        \U1/aes_core/SB3/n2469 ), .Y(\U1/aes_core/SB3/n2411 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U887  ( .A(\U1/aes_core/SB3/n2411 ), .Y(
        \U1/aes_core/SB3/n2145 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U886  ( .A(\U1/aes_core/SB3/n2402 ), .B(
        \U1/aes_core/SB3/n2475 ), .Y(\U1/aes_core/SB3/n2258 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U885  ( .A(\U1/aes_core/SB3/n2480 ), .B(
        \U1/aes_core/SB3/n2478 ), .Y(\U1/aes_core/SB3/n2436 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U883  ( .A(\U1/aes_core/SB3/n2451 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2268 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U881  ( .A0(\U1/aes_core/SB3/n2410 ), 
        .A1(\U1/aes_core/SB3/n2146 ), .B0(\U1/aes_core/SB3/n2387 ), .B1(
        \U1/aes_core/SB3/n2145 ), .C0(\U1/aes_core/SB3/n2144 ), .Y(
        \U1/aes_core/SB3/n2147 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U880  ( .AN(\U1/aes_core/SB3/n2150 ), 
        .B(\U1/aes_core/SB3/n2149 ), .C(\U1/aes_core/SB3/n2148 ), .D(
        \U1/aes_core/SB3/n2147 ), .Y(\U1/aes_core/sb3 [16]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U879  ( .A(\U1/aes_core/SB3/n2423 ), .B(
        \U1/aes_core/SB3/n2215 ), .Y(\U1/aes_core/SB3/n2275 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U878  ( .A(\U1/aes_core/SB3/n2370 ), .B(
        \U1/aes_core/SB3/n2420 ), .Y(\U1/aes_core/SB3/n2235 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U877  ( .A(\U1/aes_core/SB3/n2387 ), .B(
        \U1/aes_core/SB3/n2498 ), .Y(\U1/aes_core/SB3/n2369 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U876  ( .A0(\U1/aes_core/SB3/n2369 ), 
        .A1(\U1/aes_core/SB3/n2423 ), .B0(\U1/aes_core/SB3/n2512 ), .Y(
        \U1/aes_core/SB3/n2155 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U875  ( .A(\U1/aes_core/SB3/n2451 ), .B(
        \U1/aes_core/SB3/n2499 ), .Y(\U1/aes_core/SB3/n2251 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U874  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2451 ), .Y(\U1/aes_core/SB3/n2375 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U873  ( .A(\U1/aes_core/SB3/n2496 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2283 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U872  ( .A(\U1/aes_core/SB3/n2251 ), .B(
        \U1/aes_core/SB3/n2375 ), .C(\U1/aes_core/SB3/n2283 ), .Y(
        \U1/aes_core/SB3/n2154 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U871  ( .A(\U1/aes_core/SB3/n2451 ), .B(
        \U1/aes_core/SB3/n2510 ), .Y(\U1/aes_core/SB3/n2310 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U870  ( .A(\U1/aes_core/SB3/n2496 ), .B(
        \U1/aes_core/SB3/n2487 ), .C(\U1/aes_core/SB3/n2508 ), .Y(
        \U1/aes_core/SB3/n2151 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U869  ( .A0(\U1/aes_core/SB3/n2310 ), 
        .A1(\U1/aes_core/SB3/n2476 ), .B0(\U1/aes_core/SB3/n2151 ), .B1(
        \U1/aes_core/SB3/n2506 ), .C0(\U1/aes_core/SB3/n2370 ), .C1(
        \U1/aes_core/SB3/n2402 ), .Y(\U1/aes_core/SB3/n2153 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U868  ( .A0(\U1/aes_core/SB3/n2477 ), 
        .A1(\U1/aes_core/SB3/n2505 ), .B0(\U1/aes_core/SB3/n2478 ), .B1(
        \U1/aes_core/SB3/n2475 ), .Y(\U1/aes_core/SB3/n2152 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U867  ( .A(\U1/aes_core/SB3/n2275 ), .B(
        \U1/aes_core/SB3/n2235 ), .C(\U1/aes_core/SB3/n2155 ), .D(
        \U1/aes_core/SB3/n2154 ), .E(\U1/aes_core/SB3/n2153 ), .F(
        \U1/aes_core/SB3/n2152 ), .Y(\U1/aes_core/SB3/n2520 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U866  ( .A(\U1/aes_core/SB3/n2351 ), .B(
        \U1/aes_core/SB3/n2311 ), .Y(\U1/aes_core/SB3/n2201 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U865  ( .A0(\U1/aes_core/SB3/n2351 ), 
        .A1(\U1/aes_core/SB3/n2441 ), .B0(\U1/aes_core/SB3/n2215 ), .Y(
        \U1/aes_core/SB3/n2162 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U864  ( .A(\U1/aes_core/SB3/n2445 ), .B(
        \U1/aes_core/SB3/n2451 ), .Y(\U1/aes_core/SB3/n2203 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U863  ( .A0(\U1/aes_core/SB3/n2308 ), 
        .A1(\U1/aes_core/SB3/n2480 ), .B0(\U1/aes_core/SB3/n2203 ), .B1(
        \U1/aes_core/SB3/n2494 ), .Y(\U1/aes_core/SB3/n2161 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U862  ( .A0(\U1/aes_core/SB3/n2295 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2464 ), .B1(
        \U1/aes_core/SB3/n2370 ), .C0(\U1/aes_core/SB3/n2478 ), .C1(
        \U1/aes_core/SB3/n2421 ), .Y(\U1/aes_core/SB3/n2160 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U861  ( .A(\U1/aes_core/SB3/n2513 ), .B(
        \U1/aes_core/SB3/n2156 ), .Y(\U1/aes_core/SB3/n2259 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U860  ( .A(\U1/aes_core/SB3/n2500 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2266 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U859  ( .A(\U1/aes_core/SB3/n2442 ), .B(
        \U1/aes_core/SB3/n2495 ), .Y(\U1/aes_core/SB3/n2276 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U858  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2510 ), .Y(\U1/aes_core/SB3/n2405 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U857  ( .AN(\U1/aes_core/SB3/n2259 ), 
        .B(\U1/aes_core/SB3/n2266 ), .C(\U1/aes_core/SB3/n2276 ), .D(
        \U1/aes_core/SB3/n2405 ), .Y(\U1/aes_core/SB3/n2159 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U856  ( .A(\U1/aes_core/SB3/n2402 ), .B(
        \U1/aes_core/SB3/n2157 ), .Y(\U1/aes_core/SB3/n2384 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U855  ( .A(\U1/aes_core/SB3/n2480 ), .B(
        \U1/aes_core/SB3/n2464 ), .Y(\U1/aes_core/SB3/n2437 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U853  ( .A(\U1/aes_core/SB3/n2200 ), .B(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2225 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U851  ( .A(\U1/aes_core/SB3/n2201 ), .B(
        \U1/aes_core/SB3/n2162 ), .C(\U1/aes_core/SB3/n2161 ), .D(
        \U1/aes_core/SB3/n2160 ), .E(\U1/aes_core/SB3/n2159 ), .F(
        \U1/aes_core/SB3/n2158 ), .Y(\U1/aes_core/SB3/n2195 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U850  ( .A(\U1/aes_core/SB3/n2418 ), .B(
        \U1/aes_core/SB3/n2215 ), .Y(\U1/aes_core/SB3/n2213 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U849  ( .A(\U1/aes_core/SB3/n2370 ), .B(
        \U1/aes_core/SB3/n2295 ), .Y(\U1/aes_core/SB3/n2450 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U848  ( .A(\U1/aes_core/SB3/n2351 ), .B(
        \U1/aes_core/SB3/n2421 ), .Y(\U1/aes_core/SB3/n2263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U847  ( .A(\U1/aes_core/SB3/n2515 ), .B(
        \U1/aes_core/SB3/n2421 ), .Y(\U1/aes_core/SB3/n2278 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U846  ( .A(\U1/aes_core/SB3/n2446 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2363 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U845  ( .A(\U1/aes_core/SB3/n2496 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2230 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U844  ( .A(\U1/aes_core/SB3/n2500 ), .B(
        \U1/aes_core/SB3/n2496 ), .Y(\U1/aes_core/SB3/n2349 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U843  ( .A(\U1/aes_core/SB3/n2410 ), .B(
        \U1/aes_core/SB3/n2467 ), .Y(\U1/aes_core/SB3/n2249 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U842  ( .A(\U1/aes_core/SB3/n2363 ), .B(
        \U1/aes_core/SB3/n2230 ), .C(\U1/aes_core/SB3/n2349 ), .D(
        \U1/aes_core/SB3/n2249 ), .Y(\U1/aes_core/SB3/n2166 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U841  ( .A(\U1/aes_core/SB3/n2515 ), .B(
        \U1/aes_core/SB3/n2311 ), .Y(\U1/aes_core/SB3/n2299 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U840  ( .A(\U1/aes_core/SB3/n2514 ), .B(
        \U1/aes_core/SB3/n2295 ), .Y(\U1/aes_core/SB3/n2424 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U839  ( .A(\U1/aes_core/SB3/n2441 ), .B(
        \U1/aes_core/SB3/n2480 ), .Y(\U1/aes_core/SB3/n2374 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U838  ( .A(\U1/aes_core/SB3/n2402 ), .B(
        \U1/aes_core/SB3/n2480 ), .Y(\U1/aes_core/SB3/n2199 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U837  ( .A0(\U1/aes_core/SB3/n2480 ), 
        .A1(\U1/aes_core/SB3/n2515 ), .B0(\U1/aes_core/SB3/n2311 ), .B1(
        \U1/aes_core/SB3/n2441 ), .Y(\U1/aes_core/SB3/n2164 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U836  ( .A0(\U1/aes_core/SB3/n2295 ), 
        .A1(\U1/aes_core/SB3/n2512 ), .B0(\U1/aes_core/SB3/n2308 ), .B1(
        \U1/aes_core/SB3/n2370 ), .Y(\U1/aes_core/SB3/n2163 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U835  ( .A(\U1/aes_core/SB3/n2299 ), .B(
        \U1/aes_core/SB3/n2424 ), .C(\U1/aes_core/SB3/n2374 ), .D(
        \U1/aes_core/SB3/n2199 ), .E(\U1/aes_core/SB3/n2164 ), .F(
        \U1/aes_core/SB3/n2163 ), .Y(\U1/aes_core/SB3/n2165 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U834  ( .A(\U1/aes_core/SB3/n2213 ), .B(
        \U1/aes_core/SB3/n2450 ), .C(\U1/aes_core/SB3/n2263 ), .D(
        \U1/aes_core/SB3/n2278 ), .E(\U1/aes_core/SB3/n2166 ), .F(
        \U1/aes_core/SB3/n2165 ), .Y(\U1/aes_core/SB3/n2184 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U833  ( .A0(\U1/aes_core/SB3/n2446 ), 
        .A1(\U1/aes_core/SB3/n2443 ), .B0(\U1/aes_core/SB3/n2499 ), .B1(
        \U1/aes_core/SB3/n2387 ), .C0(\U1/aes_core/SB3/n2184 ), .Y(
        \U1/aes_core/SB3/n2167 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U832  ( .A(\U1/aes_core/SB3/n2167 ), .Y(
        \U1/aes_core/SB3/n2174 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U831  ( .A(\U1/aes_core/SB3/n2478 ), .B(
        \U1/aes_core/SB3/n2441 ), .Y(\U1/aes_core/SB3/n2468 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U830  ( .A0(\U1/aes_core/SB3/n2445 ), 
        .A1(\U1/aes_core/SB3/n2468 ), .B0(\U1/aes_core/SB3/n2500 ), .Y(
        \U1/aes_core/SB3/n2170 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U829  ( .A0(\U1/aes_core/SB3/n2410 ), 
        .A1(\U1/aes_core/SB3/n2489 ), .B0(\U1/aes_core/SB3/n2452 ), .Y(
        \U1/aes_core/SB3/n2169 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U828  ( .A0(\U1/aes_core/SB3/n2409 ), 
        .A1(\U1/aes_core/SB3/n2451 ), .B0(\U1/aes_core/SB3/n2495 ), .Y(
        \U1/aes_core/SB3/n2168 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U827  ( .A(\U1/aes_core/SB3/n2442 ), .B(
        \U1/aes_core/SB3/n2488 ), .Y(\U1/aes_core/SB3/n2242 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U826  ( .A(\U1/aes_core/SB3/n2170 ), .B(
        \U1/aes_core/SB3/n2169 ), .C(\U1/aes_core/SB3/n2168 ), .D(
        \U1/aes_core/SB3/n2242 ), .Y(\U1/aes_core/SB3/n2173 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U825  ( .A(\U1/aes_core/SB3/n2487 ), .B(
        \U1/aes_core/SB3/n2403 ), .Y(\U1/aes_core/SB3/n2457 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB3/U824  ( .A(\U1/aes_core/SB3/n2457 ), .B(
        \U1/aes_core/SB3/n2477 ), .C(\U1/aes_core/SB3/n2464 ), .Y(
        \U1/aes_core/SB3/n2171 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U823  ( .A0(\U1/aes_core/SB3/n2441 ), 
        .A1(\U1/aes_core/SB3/n2514 ), .B0(\U1/aes_core/SB3/n2171 ), .B1(
        \U1/aes_core/SB3/n2475 ), .C0(\U1/aes_core/SB3/n2513 ), .C1(
        \U1/aes_core/SB3/n2505 ), .Y(\U1/aes_core/SB3/n2172 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U822  ( .A(\U1/aes_core/SB3/n2520 ), .B(
        \U1/aes_core/SB3/n2195 ), .C(\U1/aes_core/SB3/n2175 ), .D(
        \U1/aes_core/SB3/n2174 ), .E(\U1/aes_core/SB3/n2173 ), .F(
        \U1/aes_core/SB3/n2172 ), .Y(\U1/aes_core/sb3 [17]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U821  ( .A0(\U1/aes_core/SB3/n2469 ), 
        .A1(\U1/aes_core/SB3/n2489 ), .B0(\U1/aes_core/SB3/n2510 ), .B1(
        \U1/aes_core/SB3/n2500 ), .Y(\U1/aes_core/SB3/n2176 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U820  ( .A0(\U1/aes_core/SB3/n2420 ), 
        .A1(\U1/aes_core/SB3/n2514 ), .B0(\U1/aes_core/SB3/n2370 ), .B1(
        \U1/aes_core/SB3/n2441 ), .C0(\U1/aes_core/SB3/n2176 ), .Y(
        \U1/aes_core/SB3/n2182 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U819  ( .A(\U1/aes_core/SB3/n2495 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2279 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U818  ( .A(\U1/aes_core/SB3/n2469 ), .B(
        \U1/aes_core/SB3/n2445 ), .Y(\U1/aes_core/SB3/n2260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U817  ( .A(\U1/aes_core/SB3/n2489 ), .B(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2228 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U816  ( .A(\U1/aes_core/SB3/n2409 ), .B(
        \U1/aes_core/SB3/n2452 ), .Y(\U1/aes_core/SB3/n2247 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U815  ( .A(\U1/aes_core/SB3/n2279 ), .B(
        \U1/aes_core/SB3/n2260 ), .C(\U1/aes_core/SB3/n2228 ), .D(
        \U1/aes_core/SB3/n2247 ), .Y(\U1/aes_core/SB3/n2181 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U814  ( .A(\U1/aes_core/SB3/n2515 ), .B(
        \U1/aes_core/SB3/n2493 ), .Y(\U1/aes_core/SB3/n2398 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U813  ( .A0(\U1/aes_core/SB3/n2446 ), 
        .A1(\U1/aes_core/SB3/n2398 ), .B0(\U1/aes_core/SB3/n2499 ), .Y(
        \U1/aes_core/SB3/n2179 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U812  ( .A0(\U1/aes_core/SB3/n2496 ), 
        .A1(\U1/aes_core/SB3/n2387 ), .B0(\U1/aes_core/SB3/n2399 ), .Y(
        \U1/aes_core/SB3/n2178 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U811  ( .A0(\U1/aes_core/SB3/n2404 ), 
        .A1(\U1/aes_core/SB3/n2444 ), .B0(\U1/aes_core/SB3/n2498 ), .Y(
        \U1/aes_core/SB3/n2177 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U810  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2496 ), .Y(\U1/aes_core/SB3/n2371 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U809  ( .A(\U1/aes_core/SB3/n2179 ), .B(
        \U1/aes_core/SB3/n2178 ), .C(\U1/aes_core/SB3/n2177 ), .D(
        \U1/aes_core/SB3/n2371 ), .Y(\U1/aes_core/SB3/n2180 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U808  ( .A(\U1/aes_core/SB3/n2185 ), .B(
        \U1/aes_core/SB3/n2184 ), .C(\U1/aes_core/SB3/n2183 ), .D(
        \U1/aes_core/SB3/n2182 ), .E(\U1/aes_core/SB3/n2181 ), .F(
        \U1/aes_core/SB3/n2180 ), .Y(\U1/aes_core/SB3/n2519 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U807  ( .A0(\U1/aes_core/SB3/n2300 ), 
        .A1(\U1/aes_core/SB3/n2500 ), .B0(\U1/aes_core/SB3/n2508 ), .B1(
        \U1/aes_core/SB3/n2443 ), .C0(\U1/aes_core/SB3/n2519 ), .Y(
        \U1/aes_core/SB3/n2186 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U806  ( .A(\U1/aes_core/SB3/n2186 ), .Y(
        \U1/aes_core/SB3/n2193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U805  ( .A(\U1/aes_core/SB3/n2452 ), .B(
        \U1/aes_core/SB3/n2214 ), .Y(\U1/aes_core/SB3/n2361 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U804  ( .A1N(\U1/aes_core/SB3/n2361 ), 
        .A0(\U1/aes_core/SB3/n2470 ), .B0(\U1/aes_core/SB3/n2442 ), .Y(
        \U1/aes_core/SB3/n2189 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U803  ( .A0(\U1/aes_core/SB3/n2410 ), 
        .A1(\U1/aes_core/SB3/n2293 ), .B0(\U1/aes_core/SB3/n2469 ), .Y(
        \U1/aes_core/SB3/n2188 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U802  ( .A0(\U1/aes_core/SB3/n2496 ), 
        .A1(\U1/aes_core/SB3/n2451 ), .B0(\U1/aes_core/SB3/n2490 ), .Y(
        \U1/aes_core/SB3/n2187 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U801  ( .A(\U1/aes_core/SB3/n2467 ), .B(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2243 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U800  ( .A(\U1/aes_core/SB3/n2189 ), .B(
        \U1/aes_core/SB3/n2188 ), .C(\U1/aes_core/SB3/n2187 ), .D(
        \U1/aes_core/SB3/n2243 ), .Y(\U1/aes_core/SB3/n2192 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U799  ( .A(\U1/aes_core/SB3/n2466 ), .B(
        \U1/aes_core/SB3/n2498 ), .Y(\U1/aes_core/SB3/n2497 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U798  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2444 ), .Y(\U1/aes_core/SB3/n2190 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U797  ( .A0(\U1/aes_core/SB3/n2497 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2190 ), .B1(
        \U1/aes_core/SB3/n2478 ), .C0(\U1/aes_core/SB3/n2421 ), .C1(
        \U1/aes_core/SB3/n2423 ), .Y(\U1/aes_core/SB3/n2191 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U796  ( .A(\U1/aes_core/SB3/n2196 ), .B(
        \U1/aes_core/SB3/n2195 ), .C(\U1/aes_core/SB3/n2194 ), .D(
        \U1/aes_core/SB3/n2193 ), .E(\U1/aes_core/SB3/n2192 ), .F(
        \U1/aes_core/SB3/n2191 ), .Y(\U1/aes_core/sb3 [18]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U795  ( .A(\U1/aes_core/SB3/n2300 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2502 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U794  ( .AN(\U1/aes_core/SB3/n2199 ), 
        .B(\U1/aes_core/SB3/n2198 ), .C(\U1/aes_core/SB3/n2197 ), .D(
        \U1/aes_core/SB3/n2502 ), .Y(\U1/aes_core/SB3/n2206 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U793  ( .A0(\U1/aes_core/SB3/n2200 ), 
        .A1(\U1/aes_core/SB3/n2469 ), .B0(\U1/aes_core/SB3/n2387 ), .Y(
        \U1/aes_core/SB3/n2202 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U790  ( .A(\U1/aes_core/SB3/n2443 ), .B(
        \U1/aes_core/SB3/n2490 ), .Y(\U1/aes_core/SB3/n2454 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U789  ( .A0(\U1/aes_core/SB3/n2308 ), 
        .A1(\U1/aes_core/SB3/n2512 ), .B0(\U1/aes_core/SB3/n2454 ), .B1(
        \U1/aes_core/SB3/n2465 ), .C0(\U1/aes_core/SB3/n2506 ), .C1(
        \U1/aes_core/SB3/n2515 ), .Y(\U1/aes_core/SB3/n2204 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U788  ( .A(\U1/aes_core/SB3/n2209 ), .B(
        \U1/aes_core/SB3/n2208 ), .C(\U1/aes_core/SB3/n2207 ), .D(
        \U1/aes_core/SB3/n2206 ), .E(\U1/aes_core/SB3/n2205 ), .F(
        \U1/aes_core/SB3/n2204 ), .Y(\U1/aes_core/SB3/n2417 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U787  ( .AN(\U1/aes_core/SB3/n2213 ), 
        .B(\U1/aes_core/SB3/n2212 ), .C(\U1/aes_core/SB3/n2211 ), .D(
        \U1/aes_core/SB3/n2210 ), .Y(\U1/aes_core/SB3/n2223 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U786  ( .A0(\U1/aes_core/SB3/n2500 ), 
        .A1(\U1/aes_core/SB3/n2410 ), .B0(\U1/aes_core/SB3/n2495 ), .B1(
        \U1/aes_core/SB3/n2409 ), .C0(\U1/aes_core/SB3/n2214 ), .C1(
        \U1/aes_core/SB3/n2510 ), .Y(\U1/aes_core/SB3/n2222 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U785  ( .A0(\U1/aes_core/SB3/n2464 ), 
        .A1(\U1/aes_core/SB3/n2370 ), .B0(\U1/aes_core/SB3/n2215 ), .B1(
        \U1/aes_core/SB3/n2308 ), .Y(\U1/aes_core/SB3/n2216 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U784  ( .A0(\U1/aes_core/SB3/n2387 ), 
        .A1(\U1/aes_core/SB3/n2404 ), .B0(\U1/aes_core/SB3/n2403 ), .B1(
        \U1/aes_core/SB3/n2467 ), .C0(\U1/aes_core/SB3/n2216 ), .Y(
        \U1/aes_core/SB3/n2221 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U783  ( .A(\U1/aes_core/SB3/n2475 ), .B(
        \U1/aes_core/SB3/n2514 ), .Y(\U1/aes_core/SB3/n2218 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U782  ( .A0(\U1/aes_core/SB3/n2300 ), 
        .A1(\U1/aes_core/SB3/n2219 ), .B0(\U1/aes_core/SB3/n2496 ), .B1(
        \U1/aes_core/SB3/n2218 ), .C0(\U1/aes_core/SB3/n2217 ), .Y(
        \U1/aes_core/SB3/n2220 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U781  ( .AN(\U1/aes_core/SB3/n2223 ), 
        .B(\U1/aes_core/SB3/n2222 ), .C(\U1/aes_core/SB3/n2221 ), .D(
        \U1/aes_core/SB3/n2220 ), .Y(\U1/aes_core/SB3/n2462 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U780  ( .A(\U1/aes_core/SB3/n2224 ), .Y(
        \U1/aes_core/SB3/n2240 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U779  ( .A0(\U1/aes_core/SB3/n2354 ), 
        .A1(\U1/aes_core/SB3/n2423 ), .B0(\U1/aes_core/SB3/n2225 ), .Y(
        \U1/aes_core/SB3/n2239 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U778  ( .A0(\U1/aes_core/SB3/n2496 ), 
        .A1(\U1/aes_core/SB3/n2495 ), .B0(\U1/aes_core/SB3/n2466 ), .B1(
        \U1/aes_core/SB3/n2226 ), .Y(\U1/aes_core/SB3/n2227 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U777  ( .A0(\U1/aes_core/SB3/n2477 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2493 ), .B1(
        \U1/aes_core/SB3/n2505 ), .C0(\U1/aes_core/SB3/n2227 ), .Y(
        \U1/aes_core/SB3/n2238 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U776  ( .A(\U1/aes_core/SB3/n2231 ), .B(
        \U1/aes_core/SB3/n2230 ), .C(\U1/aes_core/SB3/n2229 ), .D(
        \U1/aes_core/SB3/n2228 ), .Y(\U1/aes_core/SB3/n2237 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U775  ( .AN(\U1/aes_core/SB3/n2235 ), 
        .B(\U1/aes_core/SB3/n2234 ), .C(\U1/aes_core/SB3/n2233 ), .D(
        \U1/aes_core/SB3/n2232 ), .Y(\U1/aes_core/SB3/n2236 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U774  ( .A(\U1/aes_core/SB3/n2241 ), .B(
        \U1/aes_core/SB3/n2240 ), .C(\U1/aes_core/SB3/n2239 ), .D(
        \U1/aes_core/SB3/n2238 ), .E(\U1/aes_core/SB3/n2237 ), .F(
        \U1/aes_core/SB3/n2236 ), .Y(\U1/aes_core/SB3/n2366 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U773  ( .A0(\U1/aes_core/SB3/n2453 ), 
        .A1(\U1/aes_core/SB3/n2370 ), .B0(\U1/aes_core/SB3/n2242 ), .Y(
        \U1/aes_core/SB3/n2257 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U772  ( .AN(\U1/aes_core/SB3/n2246 ), 
        .B(\U1/aes_core/SB3/n2245 ), .C(\U1/aes_core/SB3/n2244 ), .D(
        \U1/aes_core/SB3/n2243 ), .Y(\U1/aes_core/SB3/n2256 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U771  ( .A(\U1/aes_core/SB3/n2487 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2501 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U770  ( .A(\U1/aes_core/SB3/n2249 ), .B(
        \U1/aes_core/SB3/n2248 ), .C(\U1/aes_core/SB3/n2247 ), .D(
        \U1/aes_core/SB3/n2501 ), .Y(\U1/aes_core/SB3/n2255 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U769  ( .A(\U1/aes_core/SB3/n2253 ), .B(
        \U1/aes_core/SB3/n2252 ), .C(\U1/aes_core/SB3/n2251 ), .D(
        \U1/aes_core/SB3/n2250 ), .Y(\U1/aes_core/SB3/n2254 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U768  ( .A(\U1/aes_core/SB3/n2259 ), .B(
        \U1/aes_core/SB3/n2258 ), .C(\U1/aes_core/SB3/n2257 ), .D(
        \U1/aes_core/SB3/n2256 ), .E(\U1/aes_core/SB3/n2255 ), .F(
        \U1/aes_core/SB3/n2254 ), .Y(\U1/aes_core/SB3/n2390 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U767  ( .AN(\U1/aes_core/SB3/n2263 ), 
        .B(\U1/aes_core/SB3/n2262 ), .C(\U1/aes_core/SB3/n2261 ), .D(
        \U1/aes_core/SB3/n2260 ), .Y(\U1/aes_core/SB3/n2272 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U766  ( .A(\U1/aes_core/SB3/n2267 ), .B(
        \U1/aes_core/SB3/n2266 ), .C(\U1/aes_core/SB3/n2265 ), .D(
        \U1/aes_core/SB3/n2264 ), .Y(\U1/aes_core/SB3/n2271 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U765  ( .A(\U1/aes_core/SB3/n2452 ), .B(
        \U1/aes_core/SB3/n2488 ), .C(\U1/aes_core/SB3/n2490 ), .Y(
        \U1/aes_core/SB3/n2269 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U764  ( .A0(\U1/aes_core/SB3/n2269 ), 
        .A1(\U1/aes_core/SB3/n2478 ), .B0(\U1/aes_core/SB3/n2308 ), .B1(
        \U1/aes_core/SB3/n2514 ), .C0(\U1/aes_core/SB3/n2268 ), .Y(
        \U1/aes_core/SB3/n2270 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U763  ( .A(\U1/aes_core/SB3/n2275 ), .B(
        \U1/aes_core/SB3/n2274 ), .C(\U1/aes_core/SB3/n2273 ), .D(
        \U1/aes_core/SB3/n2272 ), .E(\U1/aes_core/SB3/n2271 ), .F(
        \U1/aes_core/SB3/n2270 ), .Y(\U1/aes_core/SB3/n2438 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U762  ( .A0(\U1/aes_core/SB3/n2308 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2276 ), .Y(
        \U1/aes_core/SB3/n2290 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U761  ( .A0(\U1/aes_core/SB3/n2442 ), 
        .A1(\U1/aes_core/SB3/n2444 ), .B0(\U1/aes_core/SB3/n2499 ), .B1(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U760  ( .A0(\U1/aes_core/SB3/n2353 ), 
        .A1(\U1/aes_core/SB3/n2441 ), .B0(\U1/aes_core/SB3/n2354 ), .B1(
        \U1/aes_core/SB3/n2418 ), .C0(\U1/aes_core/SB3/n2277 ), .Y(
        \U1/aes_core/SB3/n2289 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U759  ( .A(\U1/aes_core/SB3/n2278 ), .Y(
        \U1/aes_core/SB3/n2281 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U758  ( .AN(\U1/aes_core/SB3/n2282 ), 
        .B(\U1/aes_core/SB3/n2281 ), .C(\U1/aes_core/SB3/n2280 ), .D(
        \U1/aes_core/SB3/n2279 ), .Y(\U1/aes_core/SB3/n2288 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U757  ( .A(\U1/aes_core/SB3/n2286 ), .B(
        \U1/aes_core/SB3/n2285 ), .C(\U1/aes_core/SB3/n2284 ), .D(
        \U1/aes_core/SB3/n2283 ), .Y(\U1/aes_core/SB3/n2287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U756  ( .A(\U1/aes_core/SB3/n2292 ), .B(
        \U1/aes_core/SB3/n2291 ), .C(\U1/aes_core/SB3/n2290 ), .D(
        \U1/aes_core/SB3/n2289 ), .E(\U1/aes_core/SB3/n2288 ), .F(
        \U1/aes_core/SB3/n2287 ), .Y(\U1/aes_core/SB3/n2397 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U755  ( .A0(\U1/aes_core/SB3/n2488 ), 
        .A1(\U1/aes_core/SB3/n2293 ), .B0(\U1/aes_core/SB3/n2498 ), .B1(
        \U1/aes_core/SB3/n2444 ), .Y(\U1/aes_core/SB3/n2294 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U754  ( .A0(\U1/aes_core/SB3/n2370 ), 
        .A1(\U1/aes_core/SB3/n2515 ), .B0(\U1/aes_core/SB3/n2295 ), .B1(
        \U1/aes_core/SB3/n2505 ), .C0(\U1/aes_core/SB3/n2294 ), .Y(
        \U1/aes_core/SB3/n2307 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U753  ( .AN(\U1/aes_core/SB3/n2299 ), 
        .B(\U1/aes_core/SB3/n2298 ), .C(\U1/aes_core/SB3/n2297 ), .D(
        \U1/aes_core/SB3/n2296 ), .Y(\U1/aes_core/SB3/n2306 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U752  ( .A0(\U1/aes_core/SB3/n2508 ), 
        .A1(\U1/aes_core/SB3/n2300 ), .B0(\U1/aes_core/SB3/n2499 ), .Y(
        \U1/aes_core/SB3/n2304 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U751  ( .A(\U1/aes_core/SB3/n2475 ), .B(
        \U1/aes_core/SB3/n2480 ), .Y(\U1/aes_core/SB3/n2301 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U750  ( .A0(\U1/aes_core/SB3/n2451 ), 
        .A1(\U1/aes_core/SB3/n2301 ), .B0(\U1/aes_core/SB3/n2452 ), .B1(
        \U1/aes_core/SB3/n2398 ), .Y(\U1/aes_core/SB3/n2302 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U749  ( .A(\U1/aes_core/SB3/n2304 ), .B(
        \U1/aes_core/SB3/n2303 ), .C(\U1/aes_core/SB3/n2302 ), .Y(
        \U1/aes_core/SB3/n2305 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U748  ( .A(\U1/aes_core/SB3/n2390 ), .B(
        \U1/aes_core/SB3/n2438 ), .C(\U1/aes_core/SB3/n2397 ), .D(
        \U1/aes_core/SB3/n2307 ), .E(\U1/aes_core/SB3/n2306 ), .F(
        \U1/aes_core/SB3/n2305 ), .Y(\U1/aes_core/SB3/n2484 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U747  ( .A(\U1/aes_core/SB3/n2417 ), .B(
        \U1/aes_core/SB3/n2462 ), .C(\U1/aes_core/SB3/n2366 ), .D(
        \U1/aes_core/SB3/n2484 ), .Y(\U1/aes_core/SB3/n2321 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U746  ( .A0(\U1/aes_core/SB3/n2464 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2308 ), .B1(
        \U1/aes_core/SB3/n2480 ), .Y(\U1/aes_core/SB3/n2309 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U745  ( .A0(\U1/aes_core/SB3/n2469 ), 
        .A1(\U1/aes_core/SB3/n2487 ), .B0(\U1/aes_core/SB3/n2500 ), .B1(
        \U1/aes_core/SB3/n2508 ), .C0(\U1/aes_core/SB3/n2309 ), .Y(
        \U1/aes_core/SB3/n2320 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U744  ( .A(\U1/aes_core/SB3/n2310 ), .Y(
        \U1/aes_core/SB3/n2313 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U743  ( .A0(\U1/aes_core/SB3/n2311 ), 
        .A1(\U1/aes_core/SB3/n2441 ), .B0(\U1/aes_core/SB3/n2369 ), .B1(
        \U1/aes_core/SB3/n2421 ), .Y(\U1/aes_core/SB3/n2312 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U742  ( .A0(\U1/aes_core/SB3/n2488 ), 
        .A1(\U1/aes_core/SB3/n2313 ), .B0(\U1/aes_core/SB3/n2470 ), .B1(
        \U1/aes_core/SB3/n2419 ), .C0(\U1/aes_core/SB3/n2312 ), .Y(
        \U1/aes_core/SB3/n2319 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U741  ( .A0(\U1/aes_core/SB3/n2510 ), 
        .A1(\U1/aes_core/SB3/n2387 ), .B0(\U1/aes_core/SB3/n2490 ), .Y(
        \U1/aes_core/SB3/n2317 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB3/U740  ( .A(\U1/aes_core/SB3/n2317 ), .B(
        \U1/aes_core/SB3/n2316 ), .C(\U1/aes_core/SB3/n2315 ), .D(
        \U1/aes_core/SB3/n2314 ), .Y(\U1/aes_core/SB3/n2318 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U739  ( .AN(\U1/aes_core/SB3/n2321 ), 
        .B(\U1/aes_core/SB3/n2320 ), .C(\U1/aes_core/SB3/n2319 ), .D(
        \U1/aes_core/SB3/n2318 ), .Y(\U1/aes_core/sb3 [19]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U738  ( .A(\U1/aes_core/SB3/n3166 ), .B(
        \U1/aes_core/SB3/n2983 ), .Y(\U1/aes_core/SB3/n3043 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U737  ( .A(\U1/aes_core/SB3/n3113 ), .B(
        \U1/aes_core/SB3/n3163 ), .Y(\U1/aes_core/SB3/n3003 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U736  ( .A(\U1/aes_core/SB3/n3130 ), .B(
        \U1/aes_core/SB3/n3241 ), .Y(\U1/aes_core/SB3/n3112 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U735  ( .A0(\U1/aes_core/SB3/n3112 ), 
        .A1(\U1/aes_core/SB3/n3166 ), .B0(\U1/aes_core/SB3/n3255 ), .Y(
        \U1/aes_core/SB3/n2326 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U734  ( .A(\U1/aes_core/SB3/n3194 ), .B(
        \U1/aes_core/SB3/n3242 ), .Y(\U1/aes_core/SB3/n3019 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U733  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3194 ), .Y(\U1/aes_core/SB3/n3118 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U732  ( .A(\U1/aes_core/SB3/n3239 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3051 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U731  ( .A(\U1/aes_core/SB3/n3019 ), .B(
        \U1/aes_core/SB3/n3118 ), .C(\U1/aes_core/SB3/n3051 ), .Y(
        \U1/aes_core/SB3/n2325 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U730  ( .A(\U1/aes_core/SB3/n3194 ), .B(
        \U1/aes_core/SB3/n3253 ), .Y(\U1/aes_core/SB3/n3078 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U729  ( .A(\U1/aes_core/SB3/n3239 ), .B(
        \U1/aes_core/SB3/n3230 ), .C(\U1/aes_core/SB3/n3251 ), .Y(
        \U1/aes_core/SB3/n2322 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U728  ( .A0(\U1/aes_core/SB3/n3078 ), 
        .A1(\U1/aes_core/SB3/n3219 ), .B0(\U1/aes_core/SB3/n2322 ), .B1(
        \U1/aes_core/SB3/n3249 ), .C0(\U1/aes_core/SB3/n3113 ), .C1(
        \U1/aes_core/SB3/n3145 ), .Y(\U1/aes_core/SB3/n2324 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U727  ( .A0(\U1/aes_core/SB3/n3220 ), 
        .A1(\U1/aes_core/SB3/n3248 ), .B0(\U1/aes_core/SB3/n3221 ), .B1(
        \U1/aes_core/SB3/n3218 ), .Y(\U1/aes_core/SB3/n2323 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U726  ( .A(\U1/aes_core/SB3/n3043 ), .B(
        \U1/aes_core/SB3/n3003 ), .C(\U1/aes_core/SB3/n2326 ), .D(
        \U1/aes_core/SB3/n2325 ), .E(\U1/aes_core/SB3/n2324 ), .F(
        \U1/aes_core/SB3/n2323 ), .Y(\U1/aes_core/SB3/n3263 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U725  ( .A(\U1/aes_core/SB3/n3094 ), .B(
        \U1/aes_core/SB3/n3079 ), .Y(\U1/aes_core/SB3/n2969 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U724  ( .A0(\U1/aes_core/SB3/n3094 ), 
        .A1(\U1/aes_core/SB3/n3184 ), .B0(\U1/aes_core/SB3/n2983 ), .Y(
        \U1/aes_core/SB3/n2333 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U723  ( .A(\U1/aes_core/SB3/n3188 ), .B(
        \U1/aes_core/SB3/n3194 ), .Y(\U1/aes_core/SB3/n2971 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U722  ( .A0(\U1/aes_core/SB3/n3076 ), 
        .A1(\U1/aes_core/SB3/n3223 ), .B0(\U1/aes_core/SB3/n2971 ), .B1(
        \U1/aes_core/SB3/n3237 ), .Y(\U1/aes_core/SB3/n2332 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U721  ( .A0(\U1/aes_core/SB3/n3063 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3207 ), .B1(
        \U1/aes_core/SB3/n3113 ), .C0(\U1/aes_core/SB3/n3221 ), .C1(
        \U1/aes_core/SB3/n3164 ), .Y(\U1/aes_core/SB3/n2331 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U720  ( .A(\U1/aes_core/SB3/n3256 ), .B(
        \U1/aes_core/SB3/n2327 ), .Y(\U1/aes_core/SB3/n3027 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U719  ( .A(\U1/aes_core/SB3/n3243 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3034 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U718  ( .A(\U1/aes_core/SB3/n3185 ), .B(
        \U1/aes_core/SB3/n3238 ), .Y(\U1/aes_core/SB3/n3044 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U717  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3253 ), .Y(\U1/aes_core/SB3/n3148 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U716  ( .AN(\U1/aes_core/SB3/n3027 ), 
        .B(\U1/aes_core/SB3/n3034 ), .C(\U1/aes_core/SB3/n3044 ), .D(
        \U1/aes_core/SB3/n3148 ), .Y(\U1/aes_core/SB3/n2330 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U715  ( .A(\U1/aes_core/SB3/n3145 ), .B(
        \U1/aes_core/SB3/n2328 ), .Y(\U1/aes_core/SB3/n3127 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U714  ( .A(\U1/aes_core/SB3/n3223 ), .B(
        \U1/aes_core/SB3/n3207 ), .Y(\U1/aes_core/SB3/n3180 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U712  ( .A(\U1/aes_core/SB3/n2968 ), .B(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n2993 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U710  ( .A(\U1/aes_core/SB3/n2969 ), .B(
        \U1/aes_core/SB3/n2333 ), .C(\U1/aes_core/SB3/n2332 ), .D(
        \U1/aes_core/SB3/n2331 ), .E(\U1/aes_core/SB3/n2330 ), .F(
        \U1/aes_core/SB3/n2329 ), .Y(\U1/aes_core/SB3/n2904 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U709  ( .A(\U1/aes_core/SB3/n3161 ), .B(
        \U1/aes_core/SB3/n2983 ), .Y(\U1/aes_core/SB3/n2981 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U708  ( .A(\U1/aes_core/SB3/n3113 ), .B(
        \U1/aes_core/SB3/n3063 ), .Y(\U1/aes_core/SB3/n3193 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U707  ( .A(\U1/aes_core/SB3/n3094 ), .B(
        \U1/aes_core/SB3/n3164 ), .Y(\U1/aes_core/SB3/n3031 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U706  ( .A(\U1/aes_core/SB3/n3258 ), .B(
        \U1/aes_core/SB3/n3164 ), .Y(\U1/aes_core/SB3/n3046 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U705  ( .A(\U1/aes_core/SB3/n3189 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n3106 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U704  ( .A(\U1/aes_core/SB3/n3239 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n2998 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U703  ( .A(\U1/aes_core/SB3/n3243 ), .B(
        \U1/aes_core/SB3/n3239 ), .Y(\U1/aes_core/SB3/n3092 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U702  ( .A(\U1/aes_core/SB3/n3153 ), .B(
        \U1/aes_core/SB3/n3210 ), .Y(\U1/aes_core/SB3/n3017 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U701  ( .A(\U1/aes_core/SB3/n3106 ), .B(
        \U1/aes_core/SB3/n2998 ), .C(\U1/aes_core/SB3/n3092 ), .D(
        \U1/aes_core/SB3/n3017 ), .Y(\U1/aes_core/SB3/n2337 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U700  ( .A(\U1/aes_core/SB3/n3258 ), .B(
        \U1/aes_core/SB3/n3079 ), .Y(\U1/aes_core/SB3/n3067 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U699  ( .A(\U1/aes_core/SB3/n3257 ), .B(
        \U1/aes_core/SB3/n3063 ), .Y(\U1/aes_core/SB3/n3167 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U698  ( .A(\U1/aes_core/SB3/n3184 ), .B(
        \U1/aes_core/SB3/n3223 ), .Y(\U1/aes_core/SB3/n3117 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U697  ( .A(\U1/aes_core/SB3/n3145 ), .B(
        \U1/aes_core/SB3/n3223 ), .Y(\U1/aes_core/SB3/n2967 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U696  ( .A0(\U1/aes_core/SB3/n3223 ), 
        .A1(\U1/aes_core/SB3/n3258 ), .B0(\U1/aes_core/SB3/n3079 ), .B1(
        \U1/aes_core/SB3/n3184 ), .Y(\U1/aes_core/SB3/n2335 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U695  ( .A0(\U1/aes_core/SB3/n3063 ), 
        .A1(\U1/aes_core/SB3/n3255 ), .B0(\U1/aes_core/SB3/n3076 ), .B1(
        \U1/aes_core/SB3/n3113 ), .Y(\U1/aes_core/SB3/n2334 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U694  ( .A(\U1/aes_core/SB3/n3067 ), .B(
        \U1/aes_core/SB3/n3167 ), .C(\U1/aes_core/SB3/n3117 ), .D(
        \U1/aes_core/SB3/n2967 ), .E(\U1/aes_core/SB3/n2335 ), .F(
        \U1/aes_core/SB3/n2334 ), .Y(\U1/aes_core/SB3/n2336 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U693  ( .A(\U1/aes_core/SB3/n2981 ), .B(
        \U1/aes_core/SB3/n3193 ), .C(\U1/aes_core/SB3/n3031 ), .D(
        \U1/aes_core/SB3/n3046 ), .E(\U1/aes_core/SB3/n2337 ), .F(
        \U1/aes_core/SB3/n2336 ), .Y(\U1/aes_core/SB3/n2893 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U692  ( .A0(\U1/aes_core/SB3/n3189 ), 
        .A1(\U1/aes_core/SB3/n3186 ), .B0(\U1/aes_core/SB3/n3242 ), .B1(
        \U1/aes_core/SB3/n3130 ), .C0(\U1/aes_core/SB3/n2893 ), .Y(
        \U1/aes_core/SB3/n2338 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U691  ( .A(\U1/aes_core/SB3/n2338 ), .Y(
        \U1/aes_core/SB3/n2345 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U690  ( .A(\U1/aes_core/SB3/n3221 ), .B(
        \U1/aes_core/SB3/n3184 ), .Y(\U1/aes_core/SB3/n3211 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U689  ( .A0(\U1/aes_core/SB3/n3188 ), 
        .A1(\U1/aes_core/SB3/n3211 ), .B0(\U1/aes_core/SB3/n3243 ), .Y(
        \U1/aes_core/SB3/n2341 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U688  ( .A0(\U1/aes_core/SB3/n3153 ), 
        .A1(\U1/aes_core/SB3/n3232 ), .B0(\U1/aes_core/SB3/n3195 ), .Y(
        \U1/aes_core/SB3/n2340 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U687  ( .A0(\U1/aes_core/SB3/n3152 ), 
        .A1(\U1/aes_core/SB3/n3194 ), .B0(\U1/aes_core/SB3/n3238 ), .Y(
        \U1/aes_core/SB3/n2339 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U686  ( .A(\U1/aes_core/SB3/n3185 ), .B(
        \U1/aes_core/SB3/n3231 ), .Y(\U1/aes_core/SB3/n3010 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U685  ( .A(\U1/aes_core/SB3/n2341 ), .B(
        \U1/aes_core/SB3/n2340 ), .C(\U1/aes_core/SB3/n2339 ), .D(
        \U1/aes_core/SB3/n3010 ), .Y(\U1/aes_core/SB3/n2344 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U684  ( .A(\U1/aes_core/SB3/n3230 ), .B(
        \U1/aes_core/SB3/n3146 ), .Y(\U1/aes_core/SB3/n3200 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB3/U683  ( .A(\U1/aes_core/SB3/n3200 ), .B(
        \U1/aes_core/SB3/n3220 ), .C(\U1/aes_core/SB3/n3207 ), .Y(
        \U1/aes_core/SB3/n2342 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U682  ( .A0(\U1/aes_core/SB3/n3184 ), 
        .A1(\U1/aes_core/SB3/n3257 ), .B0(\U1/aes_core/SB3/n2342 ), .B1(
        \U1/aes_core/SB3/n3218 ), .C0(\U1/aes_core/SB3/n3256 ), .C1(
        \U1/aes_core/SB3/n3248 ), .Y(\U1/aes_core/SB3/n2343 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U681  ( .A(\U1/aes_core/SB3/n3263 ), .B(
        \U1/aes_core/SB3/n2904 ), .C(\U1/aes_core/SB3/n2346 ), .D(
        \U1/aes_core/SB3/n2345 ), .E(\U1/aes_core/SB3/n2344 ), .F(
        \U1/aes_core/SB3/n2343 ), .Y(\U1/aes_core/sb3 [1]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U680  ( .A0(\U1/aes_core/SB3/n2361 ), 
        .A1(\U1/aes_core/SB3/n2476 ), .B0(\U1/aes_core/SB3/n2420 ), .Y(
        \U1/aes_core/SB3/n2358 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U679  ( .A(\U1/aes_core/SB3/n2349 ), .B(
        \U1/aes_core/SB3/n2348 ), .C(\U1/aes_core/SB3/n2347 ), .Y(
        \U1/aes_core/SB3/n2357 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U678  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2499 ), .Y(\U1/aes_core/SB3/n2352 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U677  ( .A(\U1/aes_core/SB3/n2470 ), .B(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2350 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U676  ( .A0(\U1/aes_core/SB3/n2352 ), 
        .A1(\U1/aes_core/SB3/n2351 ), .B0(\U1/aes_core/SB3/n2350 ), .B1(
        \U1/aes_core/SB3/n2493 ), .C0(\U1/aes_core/SB3/n2476 ), .C1(
        \U1/aes_core/SB3/n2402 ), .Y(\U1/aes_core/SB3/n2356 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U675  ( .A0(\U1/aes_core/SB3/n2453 ), 
        .A1(\U1/aes_core/SB3/n2354 ), .B0(\U1/aes_core/SB3/n2515 ), .B1(
        \U1/aes_core/SB3/n2505 ), .C0(\U1/aes_core/SB3/n2478 ), .C1(
        \U1/aes_core/SB3/n2353 ), .Y(\U1/aes_core/SB3/n2355 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U674  ( .A(\U1/aes_core/SB3/n2360 ), .B(
        \U1/aes_core/SB3/n2359 ), .C(\U1/aes_core/SB3/n2358 ), .D(
        \U1/aes_core/SB3/n2357 ), .E(\U1/aes_core/SB3/n2356 ), .F(
        \U1/aes_core/SB3/n2355 ), .Y(\U1/aes_core/SB3/n2485 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U673  ( .A0(\U1/aes_core/SB3/n2361 ), 
        .A1(\U1/aes_core/SB3/n2370 ), .B0(\U1/aes_core/SB3/n2441 ), .Y(
        \U1/aes_core/SB3/n2396 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB3/U672  ( .A0(\U1/aes_core/SB3/n2465 ), 
        .A1(\U1/aes_core/SB3/n2478 ), .A2(\U1/aes_core/SB3/n2418 ), .B0(
        \U1/aes_core/SB3/n2494 ), .Y(\U1/aes_core/SB3/n2395 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U671  ( .A(\U1/aes_core/SB3/n2365 ), .B(
        \U1/aes_core/SB3/n2364 ), .C(\U1/aes_core/SB3/n2363 ), .D(
        \U1/aes_core/SB3/n2362 ), .Y(\U1/aes_core/SB3/n2392 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U670  ( .A(\U1/aes_core/SB3/n2366 ), .Y(
        \U1/aes_core/SB3/n2389 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U669  ( .A(\U1/aes_core/SB3/n2367 ), .Y(
        \U1/aes_core/SB3/n2383 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB3/U668  ( .A0(\U1/aes_core/SB3/n2369 ), 
        .A1(\U1/aes_core/SB3/n2506 ), .B0N(\U1/aes_core/SB3/n2368 ), .Y(
        \U1/aes_core/SB3/n2382 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U667  ( .A0(\U1/aes_core/SB3/n2513 ), 
        .A1(\U1/aes_core/SB3/n2370 ), .B0(\U1/aes_core/SB3/n2420 ), .B1(
        \U1/aes_core/SB3/n2480 ), .C0(\U1/aes_core/SB3/n2494 ), .C1(
        \U1/aes_core/SB3/n2515 ), .Y(\U1/aes_core/SB3/n2381 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U666  ( .AN(\U1/aes_core/SB3/n2374 ), 
        .B(\U1/aes_core/SB3/n2373 ), .C(\U1/aes_core/SB3/n2372 ), .D(
        \U1/aes_core/SB3/n2371 ), .Y(\U1/aes_core/SB3/n2380 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U665  ( .A(\U1/aes_core/SB3/n2378 ), .B(
        \U1/aes_core/SB3/n2377 ), .C(\U1/aes_core/SB3/n2376 ), .D(
        \U1/aes_core/SB3/n2375 ), .Y(\U1/aes_core/SB3/n2379 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U664  ( .A(\U1/aes_core/SB3/n2384 ), .B(
        \U1/aes_core/SB3/n2383 ), .C(\U1/aes_core/SB3/n2382 ), .D(
        \U1/aes_core/SB3/n2381 ), .E(\U1/aes_core/SB3/n2380 ), .F(
        \U1/aes_core/SB3/n2379 ), .Y(\U1/aes_core/SB3/n2385 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U663  ( .A(\U1/aes_core/SB3/n2385 ), .Y(
        \U1/aes_core/SB3/n2463 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U662  ( .A0(\U1/aes_core/SB3/n2453 ), 
        .A1(\U1/aes_core/SB3/n2475 ), .B0(\U1/aes_core/SB3/n2515 ), .B1(
        \U1/aes_core/SB3/n2514 ), .Y(\U1/aes_core/SB3/n2386 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U661  ( .A0(\U1/aes_core/SB3/n2443 ), 
        .A1(\U1/aes_core/SB3/n2387 ), .B0(\U1/aes_core/SB3/n2467 ), .B1(
        \U1/aes_core/SB3/n2489 ), .C0(\U1/aes_core/SB3/n2386 ), .Y(
        \U1/aes_core/SB3/n2388 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U660  ( .AN(\U1/aes_core/SB3/n2390 ), 
        .B(\U1/aes_core/SB3/n2389 ), .C(\U1/aes_core/SB3/n2463 ), .D(
        \U1/aes_core/SB3/n2388 ), .Y(\U1/aes_core/SB3/n2391 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U659  ( .A(\U1/aes_core/SB3/n2396 ), .B(
        \U1/aes_core/SB3/n2395 ), .C(\U1/aes_core/SB3/n2394 ), .D(
        \U1/aes_core/SB3/n2393 ), .E(\U1/aes_core/SB3/n2392 ), .F(
        \U1/aes_core/SB3/n2391 ), .Y(\U1/aes_core/SB3/n2461 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U658  ( .A(\U1/aes_core/SB3/n2397 ), .Y(
        \U1/aes_core/SB3/n2401 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U657  ( .A0(\U1/aes_core/SB3/n2399 ), 
        .A1(\U1/aes_core/SB3/n2398 ), .B0(\U1/aes_core/SB3/n2445 ), .B1(
        \U1/aes_core/SB3/n2404 ), .Y(\U1/aes_core/SB3/n2400 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U656  ( .A0(\U1/aes_core/SB3/n2494 ), 
        .A1(\U1/aes_core/SB3/n2402 ), .B0(\U1/aes_core/SB3/n2401 ), .C0(
        \U1/aes_core/SB3/n2400 ), .Y(\U1/aes_core/SB3/n2416 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U655  ( .A0(\U1/aes_core/SB3/n2403 ), 
        .A1(\U1/aes_core/SB3/n2466 ), .B0(\U1/aes_core/SB3/n2495 ), .Y(
        \U1/aes_core/SB3/n2408 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U654  ( .A0(\U1/aes_core/SB3/n2404 ), 
        .A1(\U1/aes_core/SB3/n2469 ), .B0(\U1/aes_core/SB3/n2498 ), .Y(
        \U1/aes_core/SB3/n2407 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U653  ( .A(\U1/aes_core/SB3/n2408 ), .B(
        \U1/aes_core/SB3/n2407 ), .C(\U1/aes_core/SB3/n2406 ), .D(
        \U1/aes_core/SB3/n2405 ), .Y(\U1/aes_core/SB3/n2415 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U652  ( .A(\U1/aes_core/SB3/n2446 ), .B(
        \U1/aes_core/SB3/n2409 ), .Y(\U1/aes_core/SB3/n2413 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U651  ( .A(\U1/aes_core/SB3/n2410 ), .B(
        \U1/aes_core/SB3/n2451 ), .Y(\U1/aes_core/SB3/n2412 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U650  ( .A0(\U1/aes_core/SB3/n2413 ), 
        .A1(\U1/aes_core/SB3/n2512 ), .B0(\U1/aes_core/SB3/n2412 ), .B1(
        \U1/aes_core/SB3/n2476 ), .C0(\U1/aes_core/SB3/n2411 ), .C1(
        \U1/aes_core/SB3/n2477 ), .Y(\U1/aes_core/SB3/n2414 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U649  ( .A(\U1/aes_core/SB3/n2485 ), .B(
        \U1/aes_core/SB3/n2461 ), .C(\U1/aes_core/SB3/n2417 ), .D(
        \U1/aes_core/SB3/n2416 ), .E(\U1/aes_core/SB3/n2415 ), .F(
        \U1/aes_core/SB3/n2414 ), .Y(\U1/aes_core/sb3 [20]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U648  ( .A1N(\U1/aes_core/SB3/n2419 ), 
        .A0(\U1/aes_core/SB3/n2418 ), .B0(\U1/aes_core/SB3/n2475 ), .Y(
        \U1/aes_core/SB3/n2435 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U647  ( .A(\U1/aes_core/SB3/n2488 ), .B(
        \U1/aes_core/SB3/n2469 ), .Y(\U1/aes_core/SB3/n2422 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U646  ( .A0(\U1/aes_core/SB3/n2512 ), 
        .A1(\U1/aes_core/SB3/n2423 ), .B0(\U1/aes_core/SB3/n2422 ), .B1(
        \U1/aes_core/SB3/n2515 ), .C0(\U1/aes_core/SB3/n2421 ), .C1(
        \U1/aes_core/SB3/n2420 ), .Y(\U1/aes_core/SB3/n2434 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U645  ( .A(\U1/aes_core/SB3/n2424 ), .Y(
        \U1/aes_core/SB3/n2427 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U644  ( .AN(\U1/aes_core/SB3/n2428 ), 
        .B(\U1/aes_core/SB3/n2427 ), .C(\U1/aes_core/SB3/n2426 ), .D(
        \U1/aes_core/SB3/n2425 ), .Y(\U1/aes_core/SB3/n2433 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U643  ( .A(\U1/aes_core/SB3/n2431 ), .B(
        \U1/aes_core/SB3/n2430 ), .C(\U1/aes_core/SB3/n2429 ), .Y(
        \U1/aes_core/SB3/n2432 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U642  ( .A(\U1/aes_core/SB3/n2437 ), .B(
        \U1/aes_core/SB3/n2436 ), .C(\U1/aes_core/SB3/n2435 ), .D(
        \U1/aes_core/SB3/n2434 ), .E(\U1/aes_core/SB3/n2433 ), .F(
        \U1/aes_core/SB3/n2432 ), .Y(\U1/aes_core/SB3/n2486 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U641  ( .A(\U1/aes_core/SB3/n2438 ), .Y(
        \U1/aes_core/SB3/n2440 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U640  ( .A0(\U1/aes_core/SB3/n2499 ), 
        .A1(\U1/aes_core/SB3/n2496 ), .B0(\U1/aes_core/SB3/n2500 ), .B1(
        \U1/aes_core/SB3/n2498 ), .Y(\U1/aes_core/SB3/n2439 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U639  ( .A0(\U1/aes_core/SB3/n2475 ), 
        .A1(\U1/aes_core/SB3/n2441 ), .B0(\U1/aes_core/SB3/n2440 ), .C0(
        \U1/aes_core/SB3/n2439 ), .Y(\U1/aes_core/SB3/n2460 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U638  ( .A0(\U1/aes_core/SB3/n2443 ), 
        .A1(\U1/aes_core/SB3/n2499 ), .B0(\U1/aes_core/SB3/n2442 ), .Y(
        \U1/aes_core/SB3/n2449 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U637  ( .A0(\U1/aes_core/SB3/n2446 ), 
        .A1(\U1/aes_core/SB3/n2445 ), .B0(\U1/aes_core/SB3/n2444 ), .Y(
        \U1/aes_core/SB3/n2448 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U636  ( .AN(\U1/aes_core/SB3/n2450 ), 
        .B(\U1/aes_core/SB3/n2449 ), .C(\U1/aes_core/SB3/n2448 ), .D(
        \U1/aes_core/SB3/n2447 ), .Y(\U1/aes_core/SB3/n2459 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U635  ( .A0(\U1/aes_core/SB3/n2495 ), 
        .A1(\U1/aes_core/SB3/n2452 ), .B0(\U1/aes_core/SB3/n2451 ), .Y(
        \U1/aes_core/SB3/n2456 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB3/U634  ( .A0(\U1/aes_core/SB3/n2477 ), .A1(
        \U1/aes_core/SB3/n2454 ), .B0(\U1/aes_core/SB3/n2514 ), .B1(
        \U1/aes_core/SB3/n2453 ), .Y(\U1/aes_core/SB3/n2455 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U633  ( .A0(\U1/aes_core/SB3/n2457 ), 
        .A1(\U1/aes_core/SB3/n2476 ), .B0(\U1/aes_core/SB3/n2456 ), .C0(
        \U1/aes_core/SB3/n2455 ), .Y(\U1/aes_core/SB3/n2458 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U632  ( .A(\U1/aes_core/SB3/n2486 ), .B(
        \U1/aes_core/SB3/n2462 ), .C(\U1/aes_core/SB3/n2461 ), .D(
        \U1/aes_core/SB3/n2460 ), .E(\U1/aes_core/SB3/n2459 ), .F(
        \U1/aes_core/SB3/n2458 ), .Y(\U1/aes_core/sb3 [21]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U631  ( .A0(\U1/aes_core/SB3/n2465 ), 
        .A1(\U1/aes_core/SB3/n2505 ), .B0(\U1/aes_core/SB3/n2464 ), .B1(
        \U1/aes_core/SB3/n2512 ), .C0(\U1/aes_core/SB3/n2463 ), .Y(
        \U1/aes_core/SB3/n2483 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U630  ( .A0(\U1/aes_core/SB3/n2466 ), 
        .A1(\U1/aes_core/SB3/n2510 ), .B0(\U1/aes_core/SB3/n2499 ), .Y(
        \U1/aes_core/SB3/n2474 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U629  ( .A0(\U1/aes_core/SB3/n2490 ), 
        .A1(\U1/aes_core/SB3/n2467 ), .B0(\U1/aes_core/SB3/n2498 ), .Y(
        \U1/aes_core/SB3/n2473 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U628  ( .A0(\U1/aes_core/SB3/n2470 ), 
        .A1(\U1/aes_core/SB3/n2469 ), .B0(\U1/aes_core/SB3/n2468 ), .Y(
        \U1/aes_core/SB3/n2472 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U627  ( .A(\U1/aes_core/SB3/n2474 ), .B(
        \U1/aes_core/SB3/n2473 ), .C(\U1/aes_core/SB3/n2472 ), .D(
        \U1/aes_core/SB3/n2471 ), .Y(\U1/aes_core/SB3/n2482 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U626  ( .A(\U1/aes_core/SB3/n2505 ), .B(
        \U1/aes_core/SB3/n2475 ), .Y(\U1/aes_core/SB3/n2507 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U625  ( .A(\U1/aes_core/SB3/n2495 ), .B(
        \U1/aes_core/SB3/n2507 ), .Y(\U1/aes_core/SB3/n2479 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U624  ( .A0(\U1/aes_core/SB3/n2493 ), 
        .A1(\U1/aes_core/SB3/n2480 ), .B0(\U1/aes_core/SB3/n2479 ), .B1(
        \U1/aes_core/SB3/n2478 ), .C0(\U1/aes_core/SB3/n2477 ), .C1(
        \U1/aes_core/SB3/n2476 ), .Y(\U1/aes_core/SB3/n2481 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U623  ( .A(\U1/aes_core/SB3/n2486 ), .B(
        \U1/aes_core/SB3/n2485 ), .C(\U1/aes_core/SB3/n2484 ), .D(
        \U1/aes_core/SB3/n2483 ), .E(\U1/aes_core/SB3/n2482 ), .F(
        \U1/aes_core/SB3/n2481 ), .Y(\U1/aes_core/sb3 [22]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U622  ( .A0(\U1/aes_core/SB3/n2490 ), 
        .A1(\U1/aes_core/SB3/n2489 ), .B0(\U1/aes_core/SB3/n2488 ), .B1(
        \U1/aes_core/SB3/n2487 ), .Y(\U1/aes_core/SB3/n2491 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U621  ( .A0(\U1/aes_core/SB3/n2494 ), 
        .A1(\U1/aes_core/SB3/n2493 ), .B0(\U1/aes_core/SB3/n2492 ), .C0(
        \U1/aes_core/SB3/n2491 ), .Y(\U1/aes_core/SB3/n2518 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U620  ( .A1N(\U1/aes_core/SB3/n2497 ), 
        .A0(\U1/aes_core/SB3/n2496 ), .B0(\U1/aes_core/SB3/n2495 ), .Y(
        \U1/aes_core/SB3/n2504 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U619  ( .A0(\U1/aes_core/SB3/n2500 ), 
        .A1(\U1/aes_core/SB3/n2499 ), .B0(\U1/aes_core/SB3/n2498 ), .Y(
        \U1/aes_core/SB3/n2503 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U618  ( .A(\U1/aes_core/SB3/n2504 ), .B(
        \U1/aes_core/SB3/n2503 ), .C(\U1/aes_core/SB3/n2502 ), .D(
        \U1/aes_core/SB3/n2501 ), .Y(\U1/aes_core/SB3/n2517 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U617  ( .A(\U1/aes_core/SB3/n2506 ), .B(
        \U1/aes_core/SB3/n2505 ), .Y(\U1/aes_core/SB3/n2509 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U616  ( .A0(\U1/aes_core/SB3/n2510 ), 
        .A1(\U1/aes_core/SB3/n2509 ), .B0(\U1/aes_core/SB3/n2508 ), .B1(
        \U1/aes_core/SB3/n2507 ), .Y(\U1/aes_core/SB3/n2511 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U615  ( .A0(\U1/aes_core/SB3/n2515 ), 
        .A1(\U1/aes_core/SB3/n2514 ), .B0(\U1/aes_core/SB3/n2513 ), .B1(
        \U1/aes_core/SB3/n2512 ), .C0(\U1/aes_core/SB3/n2511 ), .Y(
        \U1/aes_core/SB3/n2516 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U614  ( .A(\U1/aes_core/SB3/n2521 ), .B(
        \U1/aes_core/SB3/n2520 ), .C(\U1/aes_core/SB3/n2519 ), .D(
        \U1/aes_core/SB3/n2518 ), .E(\U1/aes_core/SB3/n2517 ), .F(
        \U1/aes_core/SB3/n2516 ), .Y(\U1/aes_core/sb3 [23]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U613  ( .A(Dout[31]), .B(Dout[30]), .Y(
        \U1/aes_core/SB3/n2540 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U612  ( .A(Dout[29]), .B(Dout[28]), .Y(
        \U1/aes_core/SB3/n2531 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U611  ( .A(\U1/aes_core/SB3/n2540 ), .B(
        \U1/aes_core/SB3/n2531 ), .Y(\U1/aes_core/SB3/n2604 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U610  ( .A(Dout[25]), .Y(
        \U1/aes_core/SB3/n2525 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U609  ( .A(Dout[24]), .Y(
        \U1/aes_core/SB3/n2522 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U608  ( .A(\U1/aes_core/SB3/n2525 ), .B(
        \U1/aes_core/SB3/n2522 ), .Y(\U1/aes_core/SB3/n2532 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U607  ( .A(Dout[27]), .B(Dout[26]), .Y(
        \U1/aes_core/SB3/n2552 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U606  ( .A(\U1/aes_core/SB3/n2532 ), .B(
        \U1/aes_core/SB3/n2552 ), .Y(\U1/aes_core/SB3/n2907 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U605  ( .A(\U1/aes_core/SB3/n2604 ), .B(
        \U1/aes_core/SB3/n2907 ), .Y(\U1/aes_core/SB3/n2693 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U604  ( .A(Dout[26]), .B(Dout[27]), .Y(
        \U1/aes_core/SB3/n2535 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U603  ( .A(\U1/aes_core/SB3/n2535 ), .B(
        \U1/aes_core/SB3/n2532 ), .Y(\U1/aes_core/SB3/n2824 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U602  ( .A(Dout[31]), .Y(
        \U1/aes_core/SB3/n2528 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U601  ( .A(\U1/aes_core/SB3/n2528 ), .B(
        Dout[30]), .Y(\U1/aes_core/SB3/n2558 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U600  ( .A(\U1/aes_core/SB3/n2558 ), .B(
        \U1/aes_core/SB3/n2531 ), .Y(\U1/aes_core/SB3/n2603 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U599  ( .A(\U1/aes_core/SB3/n2824 ), .B(
        \U1/aes_core/SB3/n2603 ), .Y(\U1/aes_core/SB3/n2790 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U598  ( .A(Dout[27]), .Y(
        \U1/aes_core/SB3/n2523 ) );
  AND2_X0P5M_A12TL \U1/aes_core/SB3/U597  ( .A(Dout[26]), .B(
        \U1/aes_core/SB3/n2523 ), .Y(\U1/aes_core/SB3/n2533 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U596  ( .A(\U1/aes_core/SB3/n2532 ), .B(
        \U1/aes_core/SB3/n2533 ), .Y(\U1/aes_core/SB3/n2755 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U595  ( .A(\U1/aes_core/SB3/n2755 ), .Y(
        \U1/aes_core/SB3/n2941 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U594  ( .A(Dout[28]), .Y(
        \U1/aes_core/SB3/n2524 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U593  ( .A(\U1/aes_core/SB3/n2524 ), .B(
        Dout[29]), .Y(\U1/aes_core/SB3/n2539 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U592  ( .A(Dout[30]), .Y(
        \U1/aes_core/SB3/n2527 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U591  ( .A(\U1/aes_core/SB3/n2527 ), .B(
        Dout[31]), .Y(\U1/aes_core/SB3/n2549 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U590  ( .A(\U1/aes_core/SB3/n2539 ), .B(
        \U1/aes_core/SB3/n2549 ), .Y(\U1/aes_core/SB3/n2776 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U589  ( .A(\U1/aes_core/SB3/n2776 ), .Y(
        \U1/aes_core/SB3/n2874 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U588  ( .A(\U1/aes_core/SB3/n2941 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2733 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U587  ( .A(\U1/aes_core/SB3/n2604 ), .Y(
        \U1/aes_core/SB3/n2910 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U586  ( .A(Dout[25]), .B(Dout[24]), .Y(
        \U1/aes_core/SB3/n2536 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U585  ( .A(\U1/aes_core/SB3/n2536 ), .B(
        \U1/aes_core/SB3/n2552 ), .Y(\U1/aes_core/SB3/n2842 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U584  ( .A(\U1/aes_core/SB3/n2842 ), .Y(
        \U1/aes_core/SB3/n2951 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U583  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2951 ), .Y(\U1/aes_core/SB3/n2847 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U582  ( .A(\U1/aes_core/SB3/n2522 ), .B(
        Dout[25]), .Y(\U1/aes_core/SB3/n2551 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U581  ( .A(\U1/aes_core/SB3/n2533 ), .B(
        \U1/aes_core/SB3/n2551 ), .Y(\U1/aes_core/SB3/n2742 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U580  ( .A(\U1/aes_core/SB3/n2742 ), .Y(
        \U1/aes_core/SB3/n2831 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U579  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2711 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U578  ( .A(\U1/aes_core/SB3/n2733 ), .B(
        \U1/aes_core/SB3/n2847 ), .C(\U1/aes_core/SB3/n2711 ), .Y(
        \U1/aes_core/SB3/n2571 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U577  ( .A(\U1/aes_core/SB3/n2531 ), .B(
        \U1/aes_core/SB3/n2549 ), .Y(\U1/aes_core/SB3/n2775 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U576  ( .A(\U1/aes_core/SB3/n2523 ), .B(
        Dout[26]), .Y(\U1/aes_core/SB3/n2542 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U575  ( .A(\U1/aes_core/SB3/n2542 ), .B(
        \U1/aes_core/SB3/n2551 ), .Y(\U1/aes_core/SB3/n2773 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U574  ( .A(\U1/aes_core/SB3/n2775 ), .B(
        \U1/aes_core/SB3/n2773 ), .Y(\U1/aes_core/SB3/n2688 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U573  ( .A(\U1/aes_core/SB3/n2603 ), .Y(
        \U1/aes_core/SB3/n2912 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U572  ( .A(Dout[29]), .Y(
        \U1/aes_core/SB3/n2526 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U571  ( .A(\U1/aes_core/SB3/n2524 ), .B(
        \U1/aes_core/SB3/n2526 ), .Y(\U1/aes_core/SB3/n2550 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U570  ( .A(\U1/aes_core/SB3/n2540 ), .B(
        \U1/aes_core/SB3/n2550 ), .Y(\U1/aes_core/SB3/n2955 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U569  ( .A(\U1/aes_core/SB3/n2955 ), .Y(
        \U1/aes_core/SB3/n2865 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U568  ( .A(\U1/aes_core/SB3/n2525 ), .B(
        Dout[24]), .Y(\U1/aes_core/SB3/n2541 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U567  ( .A(\U1/aes_core/SB3/n2541 ), .B(
        \U1/aes_core/SB3/n2552 ), .Y(\U1/aes_core/SB3/n2920 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U566  ( .A(\U1/aes_core/SB3/n2920 ), .Y(
        \U1/aes_core/SB3/n2747 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U565  ( .A0(\U1/aes_core/SB3/n2912 ), 
        .A1(\U1/aes_core/SB3/n2865 ), .B0(\U1/aes_core/SB3/n2747 ), .Y(
        \U1/aes_core/SB3/n2530 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U564  ( .A(\U1/aes_core/SB3/n2536 ), .B(
        \U1/aes_core/SB3/n2533 ), .Y(\U1/aes_core/SB3/n2908 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U563  ( .A(\U1/aes_core/SB3/n2908 ), .Y(
        \U1/aes_core/SB3/n2873 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U562  ( .A(\U1/aes_core/SB3/n2526 ), .B(
        Dout[28]), .Y(\U1/aes_core/SB3/n2557 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U561  ( .A(\U1/aes_core/SB3/n2549 ), .B(
        \U1/aes_core/SB3/n2557 ), .Y(\U1/aes_core/SB3/n2948 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U560  ( .A(\U1/aes_core/SB3/n2775 ), .B(
        \U1/aes_core/SB3/n2948 ), .Y(\U1/aes_core/SB3/n2666 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U559  ( .A(\U1/aes_core/SB3/n2528 ), .B(
        \U1/aes_core/SB3/n2527 ), .Y(\U1/aes_core/SB3/n2548 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U558  ( .A(\U1/aes_core/SB3/n2539 ), .B(
        \U1/aes_core/SB3/n2548 ), .Y(\U1/aes_core/SB3/n2923 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U557  ( .A(\U1/aes_core/SB3/n2923 ), .Y(
        \U1/aes_core/SB3/n2647 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U556  ( .A0(\U1/aes_core/SB3/n2873 ), 
        .A1(\U1/aes_core/SB3/n2666 ), .B0(\U1/aes_core/SB3/n2647 ), .B1(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2529 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U555  ( .AN(\U1/aes_core/SB3/n2688 ), 
        .B(\U1/aes_core/SB3/n2530 ), .C(\U1/aes_core/SB3/n2529 ), .Y(
        \U1/aes_core/SB3/n2570 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U554  ( .A(\U1/aes_core/SB3/n2531 ), .B(
        \U1/aes_core/SB3/n2548 ), .Y(\U1/aes_core/SB3/n2792 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U553  ( .A(\U1/aes_core/SB3/n2535 ), .B(
        \U1/aes_core/SB3/n2536 ), .Y(\U1/aes_core/SB3/n2958 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U552  ( .A(\U1/aes_core/SB3/n2558 ), .B(
        \U1/aes_core/SB3/n2539 ), .Y(\U1/aes_core/SB3/n2843 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U551  ( .A(\U1/aes_core/SB3/n2535 ), .B(
        \U1/aes_core/SB3/n2541 ), .Y(\U1/aes_core/SB3/n2840 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U550  ( .A(\U1/aes_core/SB3/n2532 ), .B(
        \U1/aes_core/SB3/n2542 ), .Y(\U1/aes_core/SB3/n2845 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U549  ( .A(\U1/aes_core/SB3/n2845 ), .Y(
        \U1/aes_core/SB3/n2825 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U548  ( .A(\U1/aes_core/SB3/n2948 ), .Y(
        \U1/aes_core/SB3/n2661 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U547  ( .A(\U1/aes_core/SB3/n2533 ), .B(
        \U1/aes_core/SB3/n2541 ), .Y(\U1/aes_core/SB3/n2863 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U546  ( .A(\U1/aes_core/SB3/n2863 ), .Y(
        \U1/aes_core/SB3/n2909 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U545  ( .A0(\U1/aes_core/SB3/n2825 ), 
        .A1(\U1/aes_core/SB3/n2910 ), .B0(\U1/aes_core/SB3/n2661 ), .B1(
        \U1/aes_core/SB3/n2909 ), .Y(\U1/aes_core/SB3/n2534 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U544  ( .A0(\U1/aes_core/SB3/n2792 ), 
        .A1(\U1/aes_core/SB3/n2958 ), .B0(\U1/aes_core/SB3/n2843 ), .B1(
        \U1/aes_core/SB3/n2840 ), .C0(\U1/aes_core/SB3/n2534 ), .Y(
        \U1/aes_core/SB3/n2569 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U543  ( .A(\U1/aes_core/SB3/n2845 ), .B(
        \U1/aes_core/SB3/n2792 ), .Y(\U1/aes_core/SB3/n2654 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U542  ( .A(\U1/aes_core/SB3/n2840 ), .B(
        \U1/aes_core/SB3/n2775 ), .Y(\U1/aes_core/SB3/n2664 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U541  ( .A(\U1/aes_core/SB3/n2664 ), .Y(
        \U1/aes_core/SB3/n2538 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U540  ( .A(\U1/aes_core/SB3/n2535 ), .B(
        \U1/aes_core/SB3/n2551 ), .Y(\U1/aes_core/SB3/n2936 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U539  ( .A(\U1/aes_core/SB3/n2936 ), .Y(
        \U1/aes_core/SB3/n2864 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U538  ( .A(\U1/aes_core/SB3/n2536 ), .B(
        \U1/aes_core/SB3/n2542 ), .Y(\U1/aes_core/SB3/n2921 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U537  ( .A(\U1/aes_core/SB3/n2921 ), .Y(
        \U1/aes_core/SB3/n2932 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U536  ( .A0(\U1/aes_core/SB3/n2864 ), 
        .A1(\U1/aes_core/SB3/n2932 ), .B0(\U1/aes_core/SB3/n2865 ), .Y(
        \U1/aes_core/SB3/n2537 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U535  ( .A(\U1/aes_core/SB3/n2540 ), .B(
        \U1/aes_core/SB3/n2557 ), .Y(\U1/aes_core/SB3/n2937 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U534  ( .A(\U1/aes_core/SB3/n2937 ), .Y(
        \U1/aes_core/SB3/n2866 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U533  ( .A(\U1/aes_core/SB3/n2866 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2681 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U532  ( .AN(\U1/aes_core/SB3/n2654 ), 
        .B(\U1/aes_core/SB3/n2538 ), .C(\U1/aes_core/SB3/n2537 ), .D(
        \U1/aes_core/SB3/n2681 ), .Y(\U1/aes_core/SB3/n2547 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U531  ( .A(\U1/aes_core/SB3/n2550 ), .B(
        \U1/aes_core/SB3/n2548 ), .Y(\U1/aes_core/SB3/n2957 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U530  ( .A(\U1/aes_core/SB3/n2540 ), .B(
        \U1/aes_core/SB3/n2539 ), .Y(\U1/aes_core/SB3/n2949 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U529  ( .A0(\U1/aes_core/SB3/n2603 ), 
        .A1(\U1/aes_core/SB3/n2755 ), .B0(\U1/aes_core/SB3/n2957 ), .B1(
        \U1/aes_core/SB3/n2845 ), .C0(\U1/aes_core/SB3/n2949 ), .C1(
        \U1/aes_core/SB3/n2863 ), .Y(\U1/aes_core/SB3/n2546 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U528  ( .A(\U1/aes_core/SB3/n2908 ), .B(
        \U1/aes_core/SB3/n2603 ), .Y(\U1/aes_core/SB3/n2739 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U527  ( .A(\U1/aes_core/SB3/n2661 ), .B(
        \U1/aes_core/SB3/n2825 ), .Y(\U1/aes_core/SB3/n2692 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U526  ( .A(\U1/aes_core/SB3/n2909 ), .B(
        \U1/aes_core/SB3/n2910 ), .Y(\U1/aes_core/SB3/n2712 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U525  ( .A(\U1/aes_core/SB3/n2843 ), .Y(
        \U1/aes_core/SB3/n2938 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U524  ( .A(\U1/aes_core/SB3/n2938 ), .B(
        \U1/aes_core/SB3/n2747 ), .Y(\U1/aes_core/SB3/n2750 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U523  ( .AN(\U1/aes_core/SB3/n2739 ), 
        .B(\U1/aes_core/SB3/n2692 ), .C(\U1/aes_core/SB3/n2712 ), .D(
        \U1/aes_core/SB3/n2750 ), .Y(\U1/aes_core/SB3/n2545 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U522  ( .A(\U1/aes_core/SB3/n2558 ), .B(
        \U1/aes_core/SB3/n2550 ), .Y(\U1/aes_core/SB3/n2662 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U521  ( .A(\U1/aes_core/SB3/n2662 ), .B(
        \U1/aes_core/SB3/n2920 ), .Y(\U1/aes_core/SB3/n2816 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U520  ( .A(\U1/aes_core/SB3/n2542 ), .B(
        \U1/aes_core/SB3/n2541 ), .Y(\U1/aes_core/SB3/n2956 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U519  ( .A(\U1/aes_core/SB3/n2923 ), .B(
        \U1/aes_core/SB3/n2956 ), .Y(\U1/aes_core/SB3/n2781 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U518  ( .A(\U1/aes_core/SB3/n2781 ), .Y(
        \U1/aes_core/SB3/n2543 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U517  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2747 ), .Y(\U1/aes_core/SB3/n2800 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U516  ( .A(\U1/aes_core/SB3/n2956 ), .Y(
        \U1/aes_core/SB3/n2939 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U515  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2939 ), .Y(\U1/aes_core/SB3/n2851 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U514  ( .AN(\U1/aes_core/SB3/n2816 ), 
        .B(\U1/aes_core/SB3/n2543 ), .C(\U1/aes_core/SB3/n2800 ), .D(
        \U1/aes_core/SB3/n2851 ), .Y(\U1/aes_core/SB3/n2544 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U513  ( .A(\U1/aes_core/SB3/n2547 ), .B(
        \U1/aes_core/SB3/n2546 ), .C(\U1/aes_core/SB3/n2545 ), .D(
        \U1/aes_core/SB3/n2544 ), .Y(\U1/aes_core/SB3/n2643 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U512  ( .A(\U1/aes_core/SB3/n2842 ), .B(
        \U1/aes_core/SB3/n2662 ), .Y(\U1/aes_core/SB3/n2850 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U511  ( .A(\U1/aes_core/SB3/n2557 ), .B(
        \U1/aes_core/SB3/n2548 ), .Y(\U1/aes_core/SB3/n2758 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U510  ( .A(\U1/aes_core/SB3/n2824 ), .B(
        \U1/aes_core/SB3/n2758 ), .Y(\U1/aes_core/SB3/n2729 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U509  ( .A(\U1/aes_core/SB3/n2957 ), .Y(
        \U1/aes_core/SB3/n2913 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U508  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2873 ), .Y(\U1/aes_core/SB3/n2678 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U507  ( .A0(\U1/aes_core/SB3/n2758 ), 
        .A1(\U1/aes_core/SB3/n2956 ), .B0(\U1/aes_core/SB3/n2678 ), .Y(
        \U1/aes_core/SB3/n2556 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U506  ( .A(\U1/aes_core/SB3/n2773 ), .Y(
        \U1/aes_core/SB3/n2868 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U505  ( .A(\U1/aes_core/SB3/n2868 ), .B(
        \U1/aes_core/SB3/n2912 ), .Y(\U1/aes_core/SB3/n2869 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U504  ( .A(\U1/aes_core/SB3/n2912 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2828 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U503  ( .A(\U1/aes_core/SB3/n2550 ), .B(
        \U1/aes_core/SB3/n2549 ), .Y(\U1/aes_core/SB3/n2919 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U502  ( .A(\U1/aes_core/SB3/n2919 ), .Y(
        \U1/aes_core/SB3/n2673 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U501  ( .A(\U1/aes_core/SB3/n2864 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2697 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U500  ( .A(\U1/aes_core/SB3/n2907 ), .Y(
        \U1/aes_core/SB3/n2867 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U499  ( .A(\U1/aes_core/SB3/n2867 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2761 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U498  ( .A(\U1/aes_core/SB3/n2869 ), .B(
        \U1/aes_core/SB3/n2828 ), .C(\U1/aes_core/SB3/n2697 ), .D(
        \U1/aes_core/SB3/n2761 ), .Y(\U1/aes_core/SB3/n2555 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U497  ( .A(\U1/aes_core/SB3/n2909 ), .B(
        \U1/aes_core/SB3/n2866 ), .Y(\U1/aes_core/SB3/n2795 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U496  ( .A(\U1/aes_core/SB3/n2951 ), .B(
        \U1/aes_core/SB3/n2866 ), .Y(\U1/aes_core/SB3/n2786 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U495  ( .A(\U1/aes_core/SB3/n2949 ), .Y(
        \U1/aes_core/SB3/n2942 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U494  ( .A(\U1/aes_core/SB3/n2825 ), .B(
        \U1/aes_core/SB3/n2942 ), .Y(\U1/aes_core/SB3/n2658 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U493  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2864 ), .Y(\U1/aes_core/SB3/n2769 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U492  ( .A(\U1/aes_core/SB3/n2795 ), .B(
        \U1/aes_core/SB3/n2786 ), .C(\U1/aes_core/SB3/n2658 ), .D(
        \U1/aes_core/SB3/n2769 ), .Y(\U1/aes_core/SB3/n2554 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U491  ( .A(\U1/aes_core/SB3/n2840 ), .Y(
        \U1/aes_core/SB3/n2809 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U490  ( .A(\U1/aes_core/SB3/n2661 ), .B(
        \U1/aes_core/SB3/n2809 ), .Y(\U1/aes_core/SB3/n2645 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U489  ( .A(\U1/aes_core/SB3/n2552 ), .B(
        \U1/aes_core/SB3/n2551 ), .Y(\U1/aes_core/SB3/n2875 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U488  ( .A(\U1/aes_core/SB3/n2875 ), .Y(
        \U1/aes_core/SB3/n2930 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U487  ( .A(\U1/aes_core/SB3/n2661 ), .B(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2709 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U486  ( .A(\U1/aes_core/SB3/n2824 ), .Y(
        \U1/aes_core/SB3/n2953 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U485  ( .A(\U1/aes_core/SB3/n2953 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2744 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U484  ( .A(\U1/aes_core/SB3/n2865 ), .B(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2914 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U483  ( .A(\U1/aes_core/SB3/n2645 ), .B(
        \U1/aes_core/SB3/n2709 ), .C(\U1/aes_core/SB3/n2744 ), .D(
        \U1/aes_core/SB3/n2914 ), .Y(\U1/aes_core/SB3/n2553 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U482  ( .A(\U1/aes_core/SB3/n2850 ), .B(
        \U1/aes_core/SB3/n2729 ), .C(\U1/aes_core/SB3/n2556 ), .D(
        \U1/aes_core/SB3/n2555 ), .E(\U1/aes_core/SB3/n2554 ), .F(
        \U1/aes_core/SB3/n2553 ), .Y(\U1/aes_core/SB3/n2632 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U481  ( .A(\U1/aes_core/SB3/n2632 ), .Y(
        \U1/aes_core/SB3/n2567 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U480  ( .A(\U1/aes_core/SB3/n2921 ), .B(
        \U1/aes_core/SB3/n2758 ), .Y(\U1/aes_core/SB3/n2655 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U479  ( .A(\U1/aes_core/SB3/n2558 ), .B(
        \U1/aes_core/SB3/n2557 ), .Y(\U1/aes_core/SB3/n2918 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U478  ( .A(\U1/aes_core/SB3/n2918 ), .B(
        \U1/aes_core/SB3/n2773 ), .Y(\U1/aes_core/SB3/n2782 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U477  ( .A(\U1/aes_core/SB3/n2782 ), .Y(
        \U1/aes_core/SB3/n2560 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U476  ( .A(\U1/aes_core/SB3/n2775 ), .Y(
        \U1/aes_core/SB3/n2943 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U475  ( .A0(\U1/aes_core/SB3/n2673 ), 
        .A1(\U1/aes_core/SB3/n2943 ), .B0(\U1/aes_core/SB3/n2930 ), .Y(
        \U1/aes_core/SB3/n2559 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U474  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2809 ), .Y(\U1/aes_core/SB3/n2680 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U473  ( .AN(\U1/aes_core/SB3/n2655 ), 
        .B(\U1/aes_core/SB3/n2560 ), .C(\U1/aes_core/SB3/n2559 ), .D(
        \U1/aes_core/SB3/n2680 ), .Y(\U1/aes_core/SB3/n2564 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U472  ( .A0(\U1/aes_core/SB3/n2907 ), 
        .A1(\U1/aes_core/SB3/n2955 ), .B0(\U1/aes_core/SB3/n2792 ), .B1(
        \U1/aes_core/SB3/n2840 ), .C0(\U1/aes_core/SB3/n2920 ), .C1(
        \U1/aes_core/SB3/n2937 ), .Y(\U1/aes_core/SB3/n2563 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U471  ( .A(\U1/aes_core/SB3/n2955 ), .B(
        \U1/aes_core/SB3/n2958 ), .Y(\U1/aes_core/SB3/n2720 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U470  ( .A(\U1/aes_core/SB3/n2943 ), .B(
        \U1/aes_core/SB3/n2864 ), .Y(\U1/aes_core/SB3/n2853 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U469  ( .A(\U1/aes_core/SB3/n2825 ), .B(
        \U1/aes_core/SB3/n2943 ), .Y(\U1/aes_core/SB3/n2787 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U468  ( .A(\U1/aes_core/SB3/n2809 ), .B(
        \U1/aes_core/SB3/n2910 ), .Y(\U1/aes_core/SB3/n2659 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U467  ( .AN(\U1/aes_core/SB3/n2720 ), 
        .B(\U1/aes_core/SB3/n2853 ), .C(\U1/aes_core/SB3/n2787 ), .D(
        \U1/aes_core/SB3/n2659 ), .Y(\U1/aes_core/SB3/n2562 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U466  ( .A(\U1/aes_core/SB3/n2953 ), .B(
        \U1/aes_core/SB3/n2938 ), .Y(\U1/aes_core/SB3/n2732 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U465  ( .A(\U1/aes_core/SB3/n2809 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2799 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U464  ( .A(\U1/aes_core/SB3/n2661 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2700 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U463  ( .A(\U1/aes_core/SB3/n2868 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2745 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U462  ( .A(\U1/aes_core/SB3/n2732 ), .B(
        \U1/aes_core/SB3/n2799 ), .C(\U1/aes_core/SB3/n2700 ), .D(
        \U1/aes_core/SB3/n2745 ), .Y(\U1/aes_core/SB3/n2561 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U461  ( .A(\U1/aes_core/SB3/n2564 ), .B(
        \U1/aes_core/SB3/n2563 ), .C(\U1/aes_core/SB3/n2562 ), .D(
        \U1/aes_core/SB3/n2561 ), .Y(\U1/aes_core/SB3/n2565 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U460  ( .A(\U1/aes_core/SB3/n2565 ), .Y(
        \U1/aes_core/SB3/n2935 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U459  ( .A(\U1/aes_core/SB3/n2951 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2566 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U458  ( .AN(\U1/aes_core/SB3/n2643 ), 
        .B(\U1/aes_core/SB3/n2567 ), .C(\U1/aes_core/SB3/n2935 ), .D(
        \U1/aes_core/SB3/n2566 ), .Y(\U1/aes_core/SB3/n2568 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U457  ( .A(\U1/aes_core/SB3/n2693 ), .B(
        \U1/aes_core/SB3/n2790 ), .C(\U1/aes_core/SB3/n2571 ), .D(
        \U1/aes_core/SB3/n2570 ), .E(\U1/aes_core/SB3/n2569 ), .F(
        \U1/aes_core/SB3/n2568 ), .Y(\U1/aes_core/SB3/n2622 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U456  ( .A(\U1/aes_core/SB3/n2936 ), .B(
        \U1/aes_core/SB3/n2603 ), .Y(\U1/aes_core/SB3/n2738 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U455  ( .A(\U1/aes_core/SB3/n2865 ), .B(
        \U1/aes_core/SB3/n2953 ), .Y(\U1/aes_core/SB3/n2789 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U454  ( .A(\U1/aes_core/SB3/n2942 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2691 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U453  ( .A(\U1/aes_core/SB3/n2662 ), .Y(
        \U1/aes_core/SB3/n2931 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U452  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2714 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U451  ( .AN(\U1/aes_core/SB3/n2738 ), 
        .B(\U1/aes_core/SB3/n2789 ), .C(\U1/aes_core/SB3/n2691 ), .D(
        \U1/aes_core/SB3/n2714 ), .Y(\U1/aes_core/SB3/n2578 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U450  ( .A(\U1/aes_core/SB3/n2923 ), .B(
        \U1/aes_core/SB3/n2773 ), .Y(\U1/aes_core/SB3/n2815 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U449  ( .A(\U1/aes_core/SB3/n2825 ), .B(
        \U1/aes_core/SB3/n2912 ), .Y(\U1/aes_core/SB3/n2671 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U448  ( .A0(\U1/aes_core/SB3/n2932 ), 
        .A1(\U1/aes_core/SB3/n2831 ), .B0(\U1/aes_core/SB3/n2661 ), .Y(
        \U1/aes_core/SB3/n2572 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U447  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2763 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U446  ( .AN(\U1/aes_core/SB3/n2815 ), 
        .B(\U1/aes_core/SB3/n2671 ), .C(\U1/aes_core/SB3/n2572 ), .D(
        \U1/aes_core/SB3/n2763 ), .Y(\U1/aes_core/SB3/n2573 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U445  ( .A(\U1/aes_core/SB3/n2573 ), .Y(
        \U1/aes_core/SB3/n2577 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U444  ( .A(\U1/aes_core/SB3/n2792 ), .Y(
        \U1/aes_core/SB3/n2933 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U443  ( .A(\U1/aes_core/SB3/n2958 ), .Y(
        \U1/aes_core/SB3/n2832 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U442  ( .A0(\U1/aes_core/SB3/n2953 ), 
        .A1(\U1/aes_core/SB3/n2866 ), .B0(\U1/aes_core/SB3/n2933 ), .B1(
        \U1/aes_core/SB3/n2747 ), .C0(\U1/aes_core/SB3/n2832 ), .C1(
        \U1/aes_core/SB3/n2931 ), .Y(\U1/aes_core/SB3/n2576 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U441  ( .A0(\U1/aes_core/SB3/n2758 ), 
        .A1(\U1/aes_core/SB3/n2936 ), .B0(\U1/aes_core/SB3/n2956 ), .B1(
        \U1/aes_core/SB3/n2957 ), .Y(\U1/aes_core/SB3/n2574 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U440  ( .A0(\U1/aes_core/SB3/n2809 ), 
        .A1(\U1/aes_core/SB3/n2647 ), .B0(\U1/aes_core/SB3/n2865 ), .B1(
        \U1/aes_core/SB3/n2909 ), .C0(\U1/aes_core/SB3/n2574 ), .Y(
        \U1/aes_core/SB3/n2575 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U439  ( .AN(\U1/aes_core/SB3/n2578 ), 
        .B(\U1/aes_core/SB3/n2577 ), .C(\U1/aes_core/SB3/n2576 ), .D(
        \U1/aes_core/SB3/n2575 ), .Y(\U1/aes_core/SB3/n2641 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U438  ( .A(\U1/aes_core/SB3/n2957 ), .B(
        \U1/aes_core/SB3/n2773 ), .Y(\U1/aes_core/SB3/n2656 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U437  ( .A0(\U1/aes_core/SB3/n2843 ), 
        .A1(\U1/aes_core/SB3/n2957 ), .B0(\U1/aes_core/SB3/n2875 ), .Y(
        \U1/aes_core/SB3/n2583 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U436  ( .A(\U1/aes_core/SB3/n2875 ), .B(
        \U1/aes_core/SB3/n2863 ), .Y(\U1/aes_core/SB3/n2740 ) );
  AO22_X0P5M_A12TL \U1/aes_core/SB3/U435  ( .A0(\U1/aes_core/SB3/n2864 ), .A1(
        \U1/aes_core/SB3/n2647 ), .B0(\U1/aes_core/SB3/n2740 ), .B1(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2582 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U434  ( .A0(\U1/aes_core/SB3/n2918 ), 
        .A1(\U1/aes_core/SB3/n2958 ), .B0(\U1/aes_core/SB3/n2662 ), .B1(
        \U1/aes_core/SB3/n2755 ), .C0(\U1/aes_core/SB3/n2920 ), .C1(
        \U1/aes_core/SB3/n2949 ), .Y(\U1/aes_core/SB3/n2581 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U433  ( .A(\U1/aes_core/SB3/n2758 ), .Y(
        \U1/aes_core/SB3/n2826 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U432  ( .A(\U1/aes_core/SB3/n2951 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2852 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U431  ( .A(\U1/aes_core/SB3/n2825 ), .B(
        \U1/aes_core/SB3/n2647 ), .Y(\U1/aes_core/SB3/n2679 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U430  ( .A(\U1/aes_core/SB3/n2661 ), .B(
        \U1/aes_core/SB3/n2868 ), .Y(\U1/aes_core/SB3/n2699 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U429  ( .A(\U1/aes_core/SB3/n2825 ), .B(
        \U1/aes_core/SB3/n2866 ), .Y(\U1/aes_core/SB3/n2798 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U428  ( .A(\U1/aes_core/SB3/n2852 ), .B(
        \U1/aes_core/SB3/n2679 ), .C(\U1/aes_core/SB3/n2699 ), .D(
        \U1/aes_core/SB3/n2798 ), .Y(\U1/aes_core/SB3/n2580 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U427  ( .A(\U1/aes_core/SB3/n2845 ), .B(
        \U1/aes_core/SB3/n2758 ), .Y(\U1/aes_core/SB3/n2721 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U426  ( .A(\U1/aes_core/SB3/n2831 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2731 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U425  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2747 ), .Y(\U1/aes_core/SB3/n2762 ) );
  NAND3B_X0P5M_A12TL \U1/aes_core/SB3/U424  ( .AN(\U1/aes_core/SB3/n2721 ), 
        .B(\U1/aes_core/SB3/n2731 ), .C(\U1/aes_core/SB3/n2762 ), .Y(
        \U1/aes_core/SB3/n2579 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U423  ( .A(\U1/aes_core/SB3/n2656 ), .B(
        \U1/aes_core/SB3/n2583 ), .C(\U1/aes_core/SB3/n2582 ), .D(
        \U1/aes_core/SB3/n2581 ), .E(\U1/aes_core/SB3/n2580 ), .F(
        \U1/aes_core/SB3/n2579 ), .Y(\U1/aes_core/SB3/n2964 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U422  ( .A0(\U1/aes_core/SB3/n2661 ), 
        .A1(\U1/aes_core/SB3/n2910 ), .B0(\U1/aes_core/SB3/n2941 ), .Y(
        \U1/aes_core/SB3/n2584 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U421  ( .A(\U1/aes_core/SB3/n2647 ), .B(
        \U1/aes_core/SB3/n2747 ), .Y(\U1/aes_core/SB3/n2784 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U420  ( .A(\U1/aes_core/SB3/n2864 ), .B(
        \U1/aes_core/SB3/n2933 ), .Y(\U1/aes_core/SB3/n2676 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U419  ( .A(\U1/aes_core/SB3/n2933 ), .B(
        \U1/aes_core/SB3/n2868 ), .Y(\U1/aes_core/SB3/n2727 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U418  ( .A(\U1/aes_core/SB3/n2584 ), .B(
        \U1/aes_core/SB3/n2784 ), .C(\U1/aes_core/SB3/n2676 ), .D(
        \U1/aes_core/SB3/n2727 ), .Y(\U1/aes_core/SB3/n2588 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U417  ( .A0(\U1/aes_core/SB3/n2936 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2662 ), .B1(
        \U1/aes_core/SB3/n2908 ), .C0(\U1/aes_core/SB3/n2937 ), .C1(
        \U1/aes_core/SB3/n2773 ), .Y(\U1/aes_core/SB3/n2587 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U416  ( .A(\U1/aes_core/SB3/n2867 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2708 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U415  ( .A(\U1/aes_core/SB3/n2866 ), .B(
        \U1/aes_core/SB3/n2939 ), .Y(\U1/aes_core/SB3/n2848 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U414  ( .A(\U1/aes_core/SB3/n2866 ), .B(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2695 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U413  ( .A(\U1/aes_core/SB3/n2942 ), .B(
        \U1/aes_core/SB3/n2932 ), .Y(\U1/aes_core/SB3/n2657 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U412  ( .A(\U1/aes_core/SB3/n2708 ), .B(
        \U1/aes_core/SB3/n2848 ), .C(\U1/aes_core/SB3/n2695 ), .D(
        \U1/aes_core/SB3/n2657 ), .Y(\U1/aes_core/SB3/n2586 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U411  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2770 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U410  ( .A(\U1/aes_core/SB3/n2951 ), .B(
        \U1/aes_core/SB3/n2912 ), .Y(\U1/aes_core/SB3/n2743 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U409  ( .A(\U1/aes_core/SB3/n2941 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2794 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U408  ( .A(\U1/aes_core/SB3/n2673 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2644 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U407  ( .A(\U1/aes_core/SB3/n2770 ), .B(
        \U1/aes_core/SB3/n2743 ), .C(\U1/aes_core/SB3/n2794 ), .D(
        \U1/aes_core/SB3/n2644 ), .Y(\U1/aes_core/SB3/n2585 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U406  ( .A(\U1/aes_core/SB3/n2588 ), .B(
        \U1/aes_core/SB3/n2587 ), .C(\U1/aes_core/SB3/n2586 ), .D(
        \U1/aes_core/SB3/n2585 ), .Y(\U1/aes_core/SB3/n2630 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U405  ( .A(\U1/aes_core/SB3/n2622 ), .B(
        \U1/aes_core/SB3/n2641 ), .C(\U1/aes_core/SB3/n2964 ), .D(
        \U1/aes_core/SB3/n2630 ), .Y(\U1/aes_core/SB3/n2597 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U404  ( .A(\U1/aes_core/SB3/n2918 ), .Y(
        \U1/aes_core/SB3/n2821 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U403  ( .A0(\U1/aes_core/SB3/n2773 ), 
        .A1(\U1/aes_core/SB3/n2604 ), .B0(\U1/aes_core/SB3/n2742 ), .B1(
        \U1/aes_core/SB3/n2949 ), .Y(\U1/aes_core/SB3/n2589 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U402  ( .A0(\U1/aes_core/SB3/n2821 ), 
        .A1(\U1/aes_core/SB3/n2873 ), .B0(\U1/aes_core/SB3/n2943 ), .B1(
        \U1/aes_core/SB3/n2951 ), .C0(\U1/aes_core/SB3/n2589 ), .Y(
        \U1/aes_core/SB3/n2596 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U401  ( .A(\U1/aes_core/SB3/n2842 ), .B(
        \U1/aes_core/SB3/n2845 ), .Y(\U1/aes_core/SB3/n2841 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U400  ( .A0(\U1/aes_core/SB3/n2776 ), 
        .A1(\U1/aes_core/SB3/n2845 ), .B0(\U1/aes_core/SB3/n2758 ), .B1(
        \U1/aes_core/SB3/n2907 ), .Y(\U1/aes_core/SB3/n2590 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U399  ( .A0(\U1/aes_core/SB3/n2673 ), 
        .A1(\U1/aes_core/SB3/n2841 ), .B0(\U1/aes_core/SB3/n2913 ), .B1(
        \U1/aes_core/SB3/n2932 ), .C0(\U1/aes_core/SB3/n2590 ), .Y(
        \U1/aes_core/SB3/n2595 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U398  ( .A(\U1/aes_core/SB3/n2937 ), .B(
        \U1/aes_core/SB3/n2775 ), .Y(\U1/aes_core/SB3/n2593 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U397  ( .A(\U1/aes_core/SB3/n2866 ), .B(
        \U1/aes_core/SB3/n2912 ), .Y(\U1/aes_core/SB3/n2833 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U396  ( .A(\U1/aes_core/SB3/n2833 ), .Y(
        \U1/aes_core/SB3/n2592 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U395  ( .A(\U1/aes_core/SB3/n2824 ), .B(
        \U1/aes_core/SB3/n2918 ), .Y(\U1/aes_core/SB3/n2705 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U394  ( .A(\U1/aes_core/SB3/n2923 ), .B(
        \U1/aes_core/SB3/n2921 ), .Y(\U1/aes_core/SB3/n2858 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U392  ( .A(\U1/aes_core/SB3/n2873 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2715 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U390  ( .A0(\U1/aes_core/SB3/n2832 ), 
        .A1(\U1/aes_core/SB3/n2593 ), .B0(\U1/aes_core/SB3/n2809 ), .B1(
        \U1/aes_core/SB3/n2592 ), .C0(\U1/aes_core/SB3/n2591 ), .Y(
        \U1/aes_core/SB3/n2594 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U389  ( .AN(\U1/aes_core/SB3/n2597 ), 
        .B(\U1/aes_core/SB3/n2596 ), .C(\U1/aes_core/SB3/n2595 ), .D(
        \U1/aes_core/SB3/n2594 ), .Y(\U1/aes_core/sb3 [24]) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U388  ( .A(\U1/aes_core/SB3/n2845 ), .B(
        \U1/aes_core/SB3/n2662 ), .Y(\U1/aes_core/SB3/n2722 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U387  ( .A(\U1/aes_core/SB3/n2792 ), .B(
        \U1/aes_core/SB3/n2842 ), .Y(\U1/aes_core/SB3/n2682 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U386  ( .A(\U1/aes_core/SB3/n2809 ), .B(
        \U1/aes_core/SB3/n2941 ), .Y(\U1/aes_core/SB3/n2791 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U385  ( .A0(\U1/aes_core/SB3/n2791 ), 
        .A1(\U1/aes_core/SB3/n2845 ), .B0(\U1/aes_core/SB3/n2955 ), .Y(
        \U1/aes_core/SB3/n2602 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U384  ( .A(\U1/aes_core/SB3/n2873 ), .B(
        \U1/aes_core/SB3/n2942 ), .Y(\U1/aes_core/SB3/n2698 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U383  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2873 ), .Y(\U1/aes_core/SB3/n2797 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U382  ( .A(\U1/aes_core/SB3/n2939 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2730 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U381  ( .A(\U1/aes_core/SB3/n2698 ), .B(
        \U1/aes_core/SB3/n2797 ), .C(\U1/aes_core/SB3/n2730 ), .Y(
        \U1/aes_core/SB3/n2601 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U380  ( .A(\U1/aes_core/SB3/n2873 ), .B(
        \U1/aes_core/SB3/n2953 ), .Y(\U1/aes_core/SB3/n2757 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U379  ( .A(\U1/aes_core/SB3/n2939 ), .B(
        \U1/aes_core/SB3/n2930 ), .C(\U1/aes_core/SB3/n2951 ), .Y(
        \U1/aes_core/SB3/n2598 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U378  ( .A0(\U1/aes_core/SB3/n2757 ), 
        .A1(\U1/aes_core/SB3/n2919 ), .B0(\U1/aes_core/SB3/n2598 ), .B1(
        \U1/aes_core/SB3/n2949 ), .C0(\U1/aes_core/SB3/n2792 ), .C1(
        \U1/aes_core/SB3/n2824 ), .Y(\U1/aes_core/SB3/n2600 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U377  ( .A0(\U1/aes_core/SB3/n2920 ), 
        .A1(\U1/aes_core/SB3/n2948 ), .B0(\U1/aes_core/SB3/n2921 ), .B1(
        \U1/aes_core/SB3/n2918 ), .Y(\U1/aes_core/SB3/n2599 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U376  ( .A(\U1/aes_core/SB3/n2722 ), .B(
        \U1/aes_core/SB3/n2682 ), .C(\U1/aes_core/SB3/n2602 ), .D(
        \U1/aes_core/SB3/n2601 ), .E(\U1/aes_core/SB3/n2600 ), .F(
        \U1/aes_core/SB3/n2599 ), .Y(\U1/aes_core/SB3/n2963 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U375  ( .A(\U1/aes_core/SB3/n2773 ), .B(
        \U1/aes_core/SB3/n2758 ), .Y(\U1/aes_core/SB3/n2648 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U374  ( .A0(\U1/aes_core/SB3/n2773 ), 
        .A1(\U1/aes_core/SB3/n2863 ), .B0(\U1/aes_core/SB3/n2662 ), .Y(
        \U1/aes_core/SB3/n2609 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U373  ( .A(\U1/aes_core/SB3/n2867 ), .B(
        \U1/aes_core/SB3/n2873 ), .Y(\U1/aes_core/SB3/n2650 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U372  ( .A0(\U1/aes_core/SB3/n2755 ), 
        .A1(\U1/aes_core/SB3/n2923 ), .B0(\U1/aes_core/SB3/n2650 ), .B1(
        \U1/aes_core/SB3/n2937 ), .Y(\U1/aes_core/SB3/n2608 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U371  ( .A0(\U1/aes_core/SB3/n2742 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2907 ), .B1(
        \U1/aes_core/SB3/n2792 ), .C0(\U1/aes_core/SB3/n2921 ), .C1(
        \U1/aes_core/SB3/n2843 ), .Y(\U1/aes_core/SB3/n2607 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U370  ( .A(\U1/aes_core/SB3/n2956 ), .B(
        \U1/aes_core/SB3/n2603 ), .Y(\U1/aes_core/SB3/n2706 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U369  ( .A(\U1/aes_core/SB3/n2943 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2713 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U368  ( .A(\U1/aes_core/SB3/n2864 ), .B(
        \U1/aes_core/SB3/n2938 ), .Y(\U1/aes_core/SB3/n2723 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U367  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2953 ), .Y(\U1/aes_core/SB3/n2827 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U366  ( .AN(\U1/aes_core/SB3/n2706 ), 
        .B(\U1/aes_core/SB3/n2713 ), .C(\U1/aes_core/SB3/n2723 ), .D(
        \U1/aes_core/SB3/n2827 ), .Y(\U1/aes_core/SB3/n2606 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U365  ( .A(\U1/aes_core/SB3/n2824 ), .B(
        \U1/aes_core/SB3/n2604 ), .Y(\U1/aes_core/SB3/n2806 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U364  ( .A(\U1/aes_core/SB3/n2923 ), .B(
        \U1/aes_core/SB3/n2907 ), .Y(\U1/aes_core/SB3/n2859 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U362  ( .A(\U1/aes_core/SB3/n2647 ), .B(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2672 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U360  ( .A(\U1/aes_core/SB3/n2648 ), .B(
        \U1/aes_core/SB3/n2609 ), .C(\U1/aes_core/SB3/n2608 ), .D(
        \U1/aes_core/SB3/n2607 ), .E(\U1/aes_core/SB3/n2606 ), .F(
        \U1/aes_core/SB3/n2605 ), .Y(\U1/aes_core/SB3/n2642 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U359  ( .A(\U1/aes_core/SB3/n2840 ), .B(
        \U1/aes_core/SB3/n2662 ), .Y(\U1/aes_core/SB3/n2660 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U358  ( .A(\U1/aes_core/SB3/n2792 ), .B(
        \U1/aes_core/SB3/n2742 ), .Y(\U1/aes_core/SB3/n2872 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U357  ( .A(\U1/aes_core/SB3/n2773 ), .B(
        \U1/aes_core/SB3/n2843 ), .Y(\U1/aes_core/SB3/n2710 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U356  ( .A(\U1/aes_core/SB3/n2958 ), .B(
        \U1/aes_core/SB3/n2843 ), .Y(\U1/aes_core/SB3/n2725 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U355  ( .A(\U1/aes_core/SB3/n2868 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2785 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U354  ( .A(\U1/aes_core/SB3/n2939 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2677 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U353  ( .A(\U1/aes_core/SB3/n2943 ), .B(
        \U1/aes_core/SB3/n2939 ), .Y(\U1/aes_core/SB3/n2771 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U352  ( .A(\U1/aes_core/SB3/n2832 ), .B(
        \U1/aes_core/SB3/n2910 ), .Y(\U1/aes_core/SB3/n2696 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U351  ( .A(\U1/aes_core/SB3/n2785 ), .B(
        \U1/aes_core/SB3/n2677 ), .C(\U1/aes_core/SB3/n2771 ), .D(
        \U1/aes_core/SB3/n2696 ), .Y(\U1/aes_core/SB3/n2613 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U350  ( .A(\U1/aes_core/SB3/n2958 ), .B(
        \U1/aes_core/SB3/n2758 ), .Y(\U1/aes_core/SB3/n2746 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U349  ( .A(\U1/aes_core/SB3/n2957 ), .B(
        \U1/aes_core/SB3/n2742 ), .Y(\U1/aes_core/SB3/n2846 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U348  ( .A(\U1/aes_core/SB3/n2863 ), .B(
        \U1/aes_core/SB3/n2923 ), .Y(\U1/aes_core/SB3/n2796 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U347  ( .A(\U1/aes_core/SB3/n2824 ), .B(
        \U1/aes_core/SB3/n2923 ), .Y(\U1/aes_core/SB3/n2646 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U346  ( .A0(\U1/aes_core/SB3/n2923 ), 
        .A1(\U1/aes_core/SB3/n2958 ), .B0(\U1/aes_core/SB3/n2758 ), .B1(
        \U1/aes_core/SB3/n2863 ), .Y(\U1/aes_core/SB3/n2611 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U345  ( .A0(\U1/aes_core/SB3/n2742 ), 
        .A1(\U1/aes_core/SB3/n2955 ), .B0(\U1/aes_core/SB3/n2755 ), .B1(
        \U1/aes_core/SB3/n2792 ), .Y(\U1/aes_core/SB3/n2610 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U344  ( .A(\U1/aes_core/SB3/n2746 ), .B(
        \U1/aes_core/SB3/n2846 ), .C(\U1/aes_core/SB3/n2796 ), .D(
        \U1/aes_core/SB3/n2646 ), .E(\U1/aes_core/SB3/n2611 ), .F(
        \U1/aes_core/SB3/n2610 ), .Y(\U1/aes_core/SB3/n2612 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U343  ( .A(\U1/aes_core/SB3/n2660 ), .B(
        \U1/aes_core/SB3/n2872 ), .C(\U1/aes_core/SB3/n2710 ), .D(
        \U1/aes_core/SB3/n2725 ), .E(\U1/aes_core/SB3/n2613 ), .F(
        \U1/aes_core/SB3/n2612 ), .Y(\U1/aes_core/SB3/n2631 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U342  ( .A0(\U1/aes_core/SB3/n2868 ), 
        .A1(\U1/aes_core/SB3/n2865 ), .B0(\U1/aes_core/SB3/n2942 ), .B1(
        \U1/aes_core/SB3/n2809 ), .C0(\U1/aes_core/SB3/n2631 ), .Y(
        \U1/aes_core/SB3/n2614 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U341  ( .A(\U1/aes_core/SB3/n2614 ), .Y(
        \U1/aes_core/SB3/n2621 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U340  ( .A(\U1/aes_core/SB3/n2921 ), .B(
        \U1/aes_core/SB3/n2863 ), .Y(\U1/aes_core/SB3/n2911 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U339  ( .A0(\U1/aes_core/SB3/n2867 ), 
        .A1(\U1/aes_core/SB3/n2911 ), .B0(\U1/aes_core/SB3/n2943 ), .Y(
        \U1/aes_core/SB3/n2617 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U338  ( .A0(\U1/aes_core/SB3/n2832 ), 
        .A1(\U1/aes_core/SB3/n2932 ), .B0(\U1/aes_core/SB3/n2874 ), .Y(
        \U1/aes_core/SB3/n2616 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U337  ( .A0(\U1/aes_core/SB3/n2831 ), 
        .A1(\U1/aes_core/SB3/n2873 ), .B0(\U1/aes_core/SB3/n2938 ), .Y(
        \U1/aes_core/SB3/n2615 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U336  ( .A(\U1/aes_core/SB3/n2864 ), .B(
        \U1/aes_core/SB3/n2931 ), .Y(\U1/aes_core/SB3/n2689 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U335  ( .A(\U1/aes_core/SB3/n2617 ), .B(
        \U1/aes_core/SB3/n2616 ), .C(\U1/aes_core/SB3/n2615 ), .D(
        \U1/aes_core/SB3/n2689 ), .Y(\U1/aes_core/SB3/n2620 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U334  ( .A(\U1/aes_core/SB3/n2930 ), .B(
        \U1/aes_core/SB3/n2825 ), .Y(\U1/aes_core/SB3/n2879 ) );
  AND3_X0P5M_A12TL \U1/aes_core/SB3/U333  ( .A(\U1/aes_core/SB3/n2879 ), .B(
        \U1/aes_core/SB3/n2920 ), .C(\U1/aes_core/SB3/n2907 ), .Y(
        \U1/aes_core/SB3/n2618 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U332  ( .A0(\U1/aes_core/SB3/n2863 ), 
        .A1(\U1/aes_core/SB3/n2957 ), .B0(\U1/aes_core/SB3/n2618 ), .B1(
        \U1/aes_core/SB3/n2918 ), .C0(\U1/aes_core/SB3/n2956 ), .C1(
        \U1/aes_core/SB3/n2948 ), .Y(\U1/aes_core/SB3/n2619 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U331  ( .A(\U1/aes_core/SB3/n2963 ), .B(
        \U1/aes_core/SB3/n2642 ), .C(\U1/aes_core/SB3/n2622 ), .D(
        \U1/aes_core/SB3/n2621 ), .E(\U1/aes_core/SB3/n2620 ), .F(
        \U1/aes_core/SB3/n2619 ), .Y(\U1/aes_core/sb3 [25]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U330  ( .A0(\U1/aes_core/SB3/n2912 ), 
        .A1(\U1/aes_core/SB3/n2932 ), .B0(\U1/aes_core/SB3/n2953 ), .B1(
        \U1/aes_core/SB3/n2943 ), .Y(\U1/aes_core/SB3/n2623 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U329  ( .A0(\U1/aes_core/SB3/n2842 ), 
        .A1(\U1/aes_core/SB3/n2957 ), .B0(\U1/aes_core/SB3/n2792 ), .B1(
        \U1/aes_core/SB3/n2863 ), .C0(\U1/aes_core/SB3/n2623 ), .Y(
        \U1/aes_core/SB3/n2629 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U328  ( .A(\U1/aes_core/SB3/n2938 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2726 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U327  ( .A(\U1/aes_core/SB3/n2912 ), .B(
        \U1/aes_core/SB3/n2867 ), .Y(\U1/aes_core/SB3/n2707 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U326  ( .A(\U1/aes_core/SB3/n2932 ), .B(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2675 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U325  ( .A(\U1/aes_core/SB3/n2831 ), .B(
        \U1/aes_core/SB3/n2874 ), .Y(\U1/aes_core/SB3/n2694 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U324  ( .A(\U1/aes_core/SB3/n2726 ), .B(
        \U1/aes_core/SB3/n2707 ), .C(\U1/aes_core/SB3/n2675 ), .D(
        \U1/aes_core/SB3/n2694 ), .Y(\U1/aes_core/SB3/n2628 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U323  ( .A(\U1/aes_core/SB3/n2958 ), .B(
        \U1/aes_core/SB3/n2936 ), .Y(\U1/aes_core/SB3/n2820 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U322  ( .A0(\U1/aes_core/SB3/n2868 ), 
        .A1(\U1/aes_core/SB3/n2820 ), .B0(\U1/aes_core/SB3/n2942 ), .Y(
        \U1/aes_core/SB3/n2626 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U321  ( .A0(\U1/aes_core/SB3/n2939 ), 
        .A1(\U1/aes_core/SB3/n2809 ), .B0(\U1/aes_core/SB3/n2821 ), .Y(
        \U1/aes_core/SB3/n2625 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U320  ( .A0(\U1/aes_core/SB3/n2826 ), 
        .A1(\U1/aes_core/SB3/n2866 ), .B0(\U1/aes_core/SB3/n2941 ), .Y(
        \U1/aes_core/SB3/n2624 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U319  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2939 ), .Y(\U1/aes_core/SB3/n2793 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U318  ( .A(\U1/aes_core/SB3/n2626 ), .B(
        \U1/aes_core/SB3/n2625 ), .C(\U1/aes_core/SB3/n2624 ), .D(
        \U1/aes_core/SB3/n2793 ), .Y(\U1/aes_core/SB3/n2627 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U317  ( .A(\U1/aes_core/SB3/n2632 ), .B(
        \U1/aes_core/SB3/n2631 ), .C(\U1/aes_core/SB3/n2630 ), .D(
        \U1/aes_core/SB3/n2629 ), .E(\U1/aes_core/SB3/n2628 ), .F(
        \U1/aes_core/SB3/n2627 ), .Y(\U1/aes_core/SB3/n2962 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U316  ( .A0(\U1/aes_core/SB3/n2747 ), 
        .A1(\U1/aes_core/SB3/n2943 ), .B0(\U1/aes_core/SB3/n2951 ), .B1(
        \U1/aes_core/SB3/n2865 ), .C0(\U1/aes_core/SB3/n2962 ), .Y(
        \U1/aes_core/SB3/n2633 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U315  ( .A(\U1/aes_core/SB3/n2633 ), .Y(
        \U1/aes_core/SB3/n2640 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U314  ( .A(\U1/aes_core/SB3/n2874 ), .B(
        \U1/aes_core/SB3/n2661 ), .Y(\U1/aes_core/SB3/n2783 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U313  ( .A1N(\U1/aes_core/SB3/n2783 ), 
        .A0(\U1/aes_core/SB3/n2913 ), .B0(\U1/aes_core/SB3/n2864 ), .Y(
        \U1/aes_core/SB3/n2636 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U312  ( .A0(\U1/aes_core/SB3/n2832 ), 
        .A1(\U1/aes_core/SB3/n2740 ), .B0(\U1/aes_core/SB3/n2912 ), .Y(
        \U1/aes_core/SB3/n2635 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U311  ( .A0(\U1/aes_core/SB3/n2939 ), 
        .A1(\U1/aes_core/SB3/n2873 ), .B0(\U1/aes_core/SB3/n2933 ), .Y(
        \U1/aes_core/SB3/n2634 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U310  ( .A(\U1/aes_core/SB3/n2910 ), .B(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2690 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U309  ( .A(\U1/aes_core/SB3/n2636 ), .B(
        \U1/aes_core/SB3/n2635 ), .C(\U1/aes_core/SB3/n2634 ), .D(
        \U1/aes_core/SB3/n2690 ), .Y(\U1/aes_core/SB3/n2639 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U308  ( .A(\U1/aes_core/SB3/n2909 ), .B(
        \U1/aes_core/SB3/n2941 ), .Y(\U1/aes_core/SB3/n2940 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U307  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2866 ), .Y(\U1/aes_core/SB3/n2637 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U306  ( .A0(\U1/aes_core/SB3/n2940 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2637 ), .B1(
        \U1/aes_core/SB3/n2921 ), .C0(\U1/aes_core/SB3/n2843 ), .C1(
        \U1/aes_core/SB3/n2845 ), .Y(\U1/aes_core/SB3/n2638 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U305  ( .A(\U1/aes_core/SB3/n2643 ), .B(
        \U1/aes_core/SB3/n2642 ), .C(\U1/aes_core/SB3/n2641 ), .D(
        \U1/aes_core/SB3/n2640 ), .E(\U1/aes_core/SB3/n2639 ), .F(
        \U1/aes_core/SB3/n2638 ), .Y(\U1/aes_core/sb3 [26]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U304  ( .A(\U1/aes_core/SB3/n2747 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2945 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U303  ( .AN(\U1/aes_core/SB3/n2646 ), 
        .B(\U1/aes_core/SB3/n2645 ), .C(\U1/aes_core/SB3/n2644 ), .D(
        \U1/aes_core/SB3/n2945 ), .Y(\U1/aes_core/SB3/n2653 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U302  ( .A0(\U1/aes_core/SB3/n2647 ), 
        .A1(\U1/aes_core/SB3/n2912 ), .B0(\U1/aes_core/SB3/n2809 ), .Y(
        \U1/aes_core/SB3/n2649 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U299  ( .A(\U1/aes_core/SB3/n2865 ), .B(
        \U1/aes_core/SB3/n2933 ), .Y(\U1/aes_core/SB3/n2876 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U298  ( .A0(\U1/aes_core/SB3/n2755 ), 
        .A1(\U1/aes_core/SB3/n2955 ), .B0(\U1/aes_core/SB3/n2876 ), .B1(
        \U1/aes_core/SB3/n2908 ), .C0(\U1/aes_core/SB3/n2949 ), .C1(
        \U1/aes_core/SB3/n2958 ), .Y(\U1/aes_core/SB3/n2651 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U297  ( .A(\U1/aes_core/SB3/n2656 ), .B(
        \U1/aes_core/SB3/n2655 ), .C(\U1/aes_core/SB3/n2654 ), .D(
        \U1/aes_core/SB3/n2653 ), .E(\U1/aes_core/SB3/n2652 ), .F(
        \U1/aes_core/SB3/n2651 ), .Y(\U1/aes_core/SB3/n2839 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U296  ( .AN(\U1/aes_core/SB3/n2660 ), 
        .B(\U1/aes_core/SB3/n2659 ), .C(\U1/aes_core/SB3/n2658 ), .D(
        \U1/aes_core/SB3/n2657 ), .Y(\U1/aes_core/SB3/n2670 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U295  ( .A0(\U1/aes_core/SB3/n2943 ), 
        .A1(\U1/aes_core/SB3/n2832 ), .B0(\U1/aes_core/SB3/n2938 ), .B1(
        \U1/aes_core/SB3/n2831 ), .C0(\U1/aes_core/SB3/n2661 ), .C1(
        \U1/aes_core/SB3/n2953 ), .Y(\U1/aes_core/SB3/n2669 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U294  ( .A0(\U1/aes_core/SB3/n2907 ), 
        .A1(\U1/aes_core/SB3/n2792 ), .B0(\U1/aes_core/SB3/n2662 ), .B1(
        \U1/aes_core/SB3/n2755 ), .Y(\U1/aes_core/SB3/n2663 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U293  ( .A0(\U1/aes_core/SB3/n2809 ), 
        .A1(\U1/aes_core/SB3/n2826 ), .B0(\U1/aes_core/SB3/n2825 ), .B1(
        \U1/aes_core/SB3/n2910 ), .C0(\U1/aes_core/SB3/n2663 ), .Y(
        \U1/aes_core/SB3/n2668 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U292  ( .A(\U1/aes_core/SB3/n2918 ), .B(
        \U1/aes_core/SB3/n2957 ), .Y(\U1/aes_core/SB3/n2665 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U291  ( .A0(\U1/aes_core/SB3/n2747 ), 
        .A1(\U1/aes_core/SB3/n2666 ), .B0(\U1/aes_core/SB3/n2939 ), .B1(
        \U1/aes_core/SB3/n2665 ), .C0(\U1/aes_core/SB3/n2664 ), .Y(
        \U1/aes_core/SB3/n2667 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U290  ( .AN(\U1/aes_core/SB3/n2670 ), 
        .B(\U1/aes_core/SB3/n2669 ), .C(\U1/aes_core/SB3/n2668 ), .D(
        \U1/aes_core/SB3/n2667 ), .Y(\U1/aes_core/SB3/n2884 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U289  ( .A(\U1/aes_core/SB3/n2671 ), .Y(
        \U1/aes_core/SB3/n2687 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U288  ( .A0(\U1/aes_core/SB3/n2776 ), 
        .A1(\U1/aes_core/SB3/n2845 ), .B0(\U1/aes_core/SB3/n2672 ), .Y(
        \U1/aes_core/SB3/n2686 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U287  ( .A0(\U1/aes_core/SB3/n2939 ), 
        .A1(\U1/aes_core/SB3/n2938 ), .B0(\U1/aes_core/SB3/n2909 ), .B1(
        \U1/aes_core/SB3/n2673 ), .Y(\U1/aes_core/SB3/n2674 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U286  ( .A0(\U1/aes_core/SB3/n2920 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2936 ), .B1(
        \U1/aes_core/SB3/n2948 ), .C0(\U1/aes_core/SB3/n2674 ), .Y(
        \U1/aes_core/SB3/n2685 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U285  ( .A(\U1/aes_core/SB3/n2678 ), .B(
        \U1/aes_core/SB3/n2677 ), .C(\U1/aes_core/SB3/n2676 ), .D(
        \U1/aes_core/SB3/n2675 ), .Y(\U1/aes_core/SB3/n2684 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U284  ( .AN(\U1/aes_core/SB3/n2682 ), 
        .B(\U1/aes_core/SB3/n2681 ), .C(\U1/aes_core/SB3/n2680 ), .D(
        \U1/aes_core/SB3/n2679 ), .Y(\U1/aes_core/SB3/n2683 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U283  ( .A(\U1/aes_core/SB3/n2688 ), .B(
        \U1/aes_core/SB3/n2687 ), .C(\U1/aes_core/SB3/n2686 ), .D(
        \U1/aes_core/SB3/n2685 ), .E(\U1/aes_core/SB3/n2684 ), .F(
        \U1/aes_core/SB3/n2683 ), .Y(\U1/aes_core/SB3/n2788 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U282  ( .A0(\U1/aes_core/SB3/n2875 ), 
        .A1(\U1/aes_core/SB3/n2792 ), .B0(\U1/aes_core/SB3/n2689 ), .Y(
        \U1/aes_core/SB3/n2704 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U281  ( .AN(\U1/aes_core/SB3/n2693 ), 
        .B(\U1/aes_core/SB3/n2692 ), .C(\U1/aes_core/SB3/n2691 ), .D(
        \U1/aes_core/SB3/n2690 ), .Y(\U1/aes_core/SB3/n2703 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U280  ( .A(\U1/aes_core/SB3/n2930 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2944 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U279  ( .A(\U1/aes_core/SB3/n2696 ), .B(
        \U1/aes_core/SB3/n2695 ), .C(\U1/aes_core/SB3/n2694 ), .D(
        \U1/aes_core/SB3/n2944 ), .Y(\U1/aes_core/SB3/n2702 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U278  ( .A(\U1/aes_core/SB3/n2700 ), .B(
        \U1/aes_core/SB3/n2699 ), .C(\U1/aes_core/SB3/n2698 ), .D(
        \U1/aes_core/SB3/n2697 ), .Y(\U1/aes_core/SB3/n2701 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U277  ( .A(\U1/aes_core/SB3/n2706 ), .B(
        \U1/aes_core/SB3/n2705 ), .C(\U1/aes_core/SB3/n2704 ), .D(
        \U1/aes_core/SB3/n2703 ), .E(\U1/aes_core/SB3/n2702 ), .F(
        \U1/aes_core/SB3/n2701 ), .Y(\U1/aes_core/SB3/n2812 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U276  ( .AN(\U1/aes_core/SB3/n2710 ), 
        .B(\U1/aes_core/SB3/n2709 ), .C(\U1/aes_core/SB3/n2708 ), .D(
        \U1/aes_core/SB3/n2707 ), .Y(\U1/aes_core/SB3/n2719 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U275  ( .A(\U1/aes_core/SB3/n2714 ), .B(
        \U1/aes_core/SB3/n2713 ), .C(\U1/aes_core/SB3/n2712 ), .D(
        \U1/aes_core/SB3/n2711 ), .Y(\U1/aes_core/SB3/n2718 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U274  ( .A(\U1/aes_core/SB3/n2874 ), .B(
        \U1/aes_core/SB3/n2931 ), .C(\U1/aes_core/SB3/n2933 ), .Y(
        \U1/aes_core/SB3/n2716 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U273  ( .A0(\U1/aes_core/SB3/n2716 ), 
        .A1(\U1/aes_core/SB3/n2921 ), .B0(\U1/aes_core/SB3/n2755 ), .B1(
        \U1/aes_core/SB3/n2957 ), .C0(\U1/aes_core/SB3/n2715 ), .Y(
        \U1/aes_core/SB3/n2717 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U272  ( .A(\U1/aes_core/SB3/n2722 ), .B(
        \U1/aes_core/SB3/n2721 ), .C(\U1/aes_core/SB3/n2720 ), .D(
        \U1/aes_core/SB3/n2719 ), .E(\U1/aes_core/SB3/n2718 ), .F(
        \U1/aes_core/SB3/n2717 ), .Y(\U1/aes_core/SB3/n2860 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U271  ( .A0(\U1/aes_core/SB3/n2755 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2723 ), .Y(
        \U1/aes_core/SB3/n2737 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U270  ( .A0(\U1/aes_core/SB3/n2864 ), 
        .A1(\U1/aes_core/SB3/n2866 ), .B0(\U1/aes_core/SB3/n2942 ), .B1(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2724 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U269  ( .A0(\U1/aes_core/SB3/n2775 ), 
        .A1(\U1/aes_core/SB3/n2863 ), .B0(\U1/aes_core/SB3/n2776 ), .B1(
        \U1/aes_core/SB3/n2840 ), .C0(\U1/aes_core/SB3/n2724 ), .Y(
        \U1/aes_core/SB3/n2736 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U268  ( .A(\U1/aes_core/SB3/n2725 ), .Y(
        \U1/aes_core/SB3/n2728 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U267  ( .AN(\U1/aes_core/SB3/n2729 ), 
        .B(\U1/aes_core/SB3/n2728 ), .C(\U1/aes_core/SB3/n2727 ), .D(
        \U1/aes_core/SB3/n2726 ), .Y(\U1/aes_core/SB3/n2735 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U266  ( .A(\U1/aes_core/SB3/n2733 ), .B(
        \U1/aes_core/SB3/n2732 ), .C(\U1/aes_core/SB3/n2731 ), .D(
        \U1/aes_core/SB3/n2730 ), .Y(\U1/aes_core/SB3/n2734 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U265  ( .A(\U1/aes_core/SB3/n2739 ), .B(
        \U1/aes_core/SB3/n2738 ), .C(\U1/aes_core/SB3/n2737 ), .D(
        \U1/aes_core/SB3/n2736 ), .E(\U1/aes_core/SB3/n2735 ), .F(
        \U1/aes_core/SB3/n2734 ), .Y(\U1/aes_core/SB3/n2819 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U264  ( .A0(\U1/aes_core/SB3/n2931 ), 
        .A1(\U1/aes_core/SB3/n2740 ), .B0(\U1/aes_core/SB3/n2941 ), .B1(
        \U1/aes_core/SB3/n2866 ), .Y(\U1/aes_core/SB3/n2741 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U263  ( .A0(\U1/aes_core/SB3/n2792 ), 
        .A1(\U1/aes_core/SB3/n2958 ), .B0(\U1/aes_core/SB3/n2742 ), .B1(
        \U1/aes_core/SB3/n2948 ), .C0(\U1/aes_core/SB3/n2741 ), .Y(
        \U1/aes_core/SB3/n2754 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U262  ( .AN(\U1/aes_core/SB3/n2746 ), 
        .B(\U1/aes_core/SB3/n2745 ), .C(\U1/aes_core/SB3/n2744 ), .D(
        \U1/aes_core/SB3/n2743 ), .Y(\U1/aes_core/SB3/n2753 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U261  ( .A0(\U1/aes_core/SB3/n2951 ), 
        .A1(\U1/aes_core/SB3/n2747 ), .B0(\U1/aes_core/SB3/n2942 ), .Y(
        \U1/aes_core/SB3/n2751 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U260  ( .A(\U1/aes_core/SB3/n2918 ), .B(
        \U1/aes_core/SB3/n2923 ), .Y(\U1/aes_core/SB3/n2748 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U259  ( .A0(\U1/aes_core/SB3/n2873 ), 
        .A1(\U1/aes_core/SB3/n2748 ), .B0(\U1/aes_core/SB3/n2874 ), .B1(
        \U1/aes_core/SB3/n2820 ), .Y(\U1/aes_core/SB3/n2749 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U258  ( .A(\U1/aes_core/SB3/n2751 ), .B(
        \U1/aes_core/SB3/n2750 ), .C(\U1/aes_core/SB3/n2749 ), .Y(
        \U1/aes_core/SB3/n2752 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U257  ( .A(\U1/aes_core/SB3/n2812 ), .B(
        \U1/aes_core/SB3/n2860 ), .C(\U1/aes_core/SB3/n2819 ), .D(
        \U1/aes_core/SB3/n2754 ), .E(\U1/aes_core/SB3/n2753 ), .F(
        \U1/aes_core/SB3/n2752 ), .Y(\U1/aes_core/SB3/n2927 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U256  ( .A(\U1/aes_core/SB3/n2839 ), .B(
        \U1/aes_core/SB3/n2884 ), .C(\U1/aes_core/SB3/n2788 ), .D(
        \U1/aes_core/SB3/n2927 ), .Y(\U1/aes_core/SB3/n2768 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U255  ( .A0(\U1/aes_core/SB3/n2907 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2755 ), .B1(
        \U1/aes_core/SB3/n2923 ), .Y(\U1/aes_core/SB3/n2756 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U254  ( .A0(\U1/aes_core/SB3/n2912 ), 
        .A1(\U1/aes_core/SB3/n2930 ), .B0(\U1/aes_core/SB3/n2943 ), .B1(
        \U1/aes_core/SB3/n2951 ), .C0(\U1/aes_core/SB3/n2756 ), .Y(
        \U1/aes_core/SB3/n2767 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U253  ( .A(\U1/aes_core/SB3/n2757 ), .Y(
        \U1/aes_core/SB3/n2760 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U252  ( .A0(\U1/aes_core/SB3/n2758 ), 
        .A1(\U1/aes_core/SB3/n2863 ), .B0(\U1/aes_core/SB3/n2791 ), .B1(
        \U1/aes_core/SB3/n2843 ), .Y(\U1/aes_core/SB3/n2759 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U251  ( .A0(\U1/aes_core/SB3/n2931 ), 
        .A1(\U1/aes_core/SB3/n2760 ), .B0(\U1/aes_core/SB3/n2913 ), .B1(
        \U1/aes_core/SB3/n2841 ), .C0(\U1/aes_core/SB3/n2759 ), .Y(
        \U1/aes_core/SB3/n2766 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U250  ( .A0(\U1/aes_core/SB3/n2953 ), 
        .A1(\U1/aes_core/SB3/n2809 ), .B0(\U1/aes_core/SB3/n2933 ), .Y(
        \U1/aes_core/SB3/n2764 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB3/U249  ( .A(\U1/aes_core/SB3/n2764 ), .B(
        \U1/aes_core/SB3/n2763 ), .C(\U1/aes_core/SB3/n2762 ), .D(
        \U1/aes_core/SB3/n2761 ), .Y(\U1/aes_core/SB3/n2765 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U248  ( .AN(\U1/aes_core/SB3/n2768 ), 
        .B(\U1/aes_core/SB3/n2767 ), .C(\U1/aes_core/SB3/n2766 ), .D(
        \U1/aes_core/SB3/n2765 ), .Y(\U1/aes_core/sb3 [27]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U247  ( .A0(\U1/aes_core/SB3/n2783 ), 
        .A1(\U1/aes_core/SB3/n2919 ), .B0(\U1/aes_core/SB3/n2842 ), .Y(
        \U1/aes_core/SB3/n2780 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U246  ( .A(\U1/aes_core/SB3/n2771 ), .B(
        \U1/aes_core/SB3/n2770 ), .C(\U1/aes_core/SB3/n2769 ), .Y(
        \U1/aes_core/SB3/n2779 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U245  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2942 ), .Y(\U1/aes_core/SB3/n2774 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U244  ( .A(\U1/aes_core/SB3/n2913 ), .B(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2772 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U243  ( .A0(\U1/aes_core/SB3/n2774 ), 
        .A1(\U1/aes_core/SB3/n2773 ), .B0(\U1/aes_core/SB3/n2772 ), .B1(
        \U1/aes_core/SB3/n2936 ), .C0(\U1/aes_core/SB3/n2919 ), .C1(
        \U1/aes_core/SB3/n2824 ), .Y(\U1/aes_core/SB3/n2778 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U242  ( .A0(\U1/aes_core/SB3/n2875 ), 
        .A1(\U1/aes_core/SB3/n2776 ), .B0(\U1/aes_core/SB3/n2958 ), .B1(
        \U1/aes_core/SB3/n2948 ), .C0(\U1/aes_core/SB3/n2921 ), .C1(
        \U1/aes_core/SB3/n2775 ), .Y(\U1/aes_core/SB3/n2777 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U241  ( .A(\U1/aes_core/SB3/n2782 ), .B(
        \U1/aes_core/SB3/n2781 ), .C(\U1/aes_core/SB3/n2780 ), .D(
        \U1/aes_core/SB3/n2779 ), .E(\U1/aes_core/SB3/n2778 ), .F(
        \U1/aes_core/SB3/n2777 ), .Y(\U1/aes_core/SB3/n2928 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U240  ( .A0(\U1/aes_core/SB3/n2783 ), 
        .A1(\U1/aes_core/SB3/n2792 ), .B0(\U1/aes_core/SB3/n2863 ), .Y(
        \U1/aes_core/SB3/n2818 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB3/U239  ( .A0(\U1/aes_core/SB3/n2908 ), 
        .A1(\U1/aes_core/SB3/n2921 ), .A2(\U1/aes_core/SB3/n2840 ), .B0(
        \U1/aes_core/SB3/n2937 ), .Y(\U1/aes_core/SB3/n2817 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U238  ( .A(\U1/aes_core/SB3/n2787 ), .B(
        \U1/aes_core/SB3/n2786 ), .C(\U1/aes_core/SB3/n2785 ), .D(
        \U1/aes_core/SB3/n2784 ), .Y(\U1/aes_core/SB3/n2814 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U237  ( .A(\U1/aes_core/SB3/n2788 ), .Y(
        \U1/aes_core/SB3/n2811 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U236  ( .A(\U1/aes_core/SB3/n2789 ), .Y(
        \U1/aes_core/SB3/n2805 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB3/U235  ( .A0(\U1/aes_core/SB3/n2791 ), 
        .A1(\U1/aes_core/SB3/n2949 ), .B0N(\U1/aes_core/SB3/n2790 ), .Y(
        \U1/aes_core/SB3/n2804 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U234  ( .A0(\U1/aes_core/SB3/n2956 ), 
        .A1(\U1/aes_core/SB3/n2792 ), .B0(\U1/aes_core/SB3/n2842 ), .B1(
        \U1/aes_core/SB3/n2923 ), .C0(\U1/aes_core/SB3/n2937 ), .C1(
        \U1/aes_core/SB3/n2958 ), .Y(\U1/aes_core/SB3/n2803 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U233  ( .AN(\U1/aes_core/SB3/n2796 ), 
        .B(\U1/aes_core/SB3/n2795 ), .C(\U1/aes_core/SB3/n2794 ), .D(
        \U1/aes_core/SB3/n2793 ), .Y(\U1/aes_core/SB3/n2802 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U232  ( .A(\U1/aes_core/SB3/n2800 ), .B(
        \U1/aes_core/SB3/n2799 ), .C(\U1/aes_core/SB3/n2798 ), .D(
        \U1/aes_core/SB3/n2797 ), .Y(\U1/aes_core/SB3/n2801 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U231  ( .A(\U1/aes_core/SB3/n2806 ), .B(
        \U1/aes_core/SB3/n2805 ), .C(\U1/aes_core/SB3/n2804 ), .D(
        \U1/aes_core/SB3/n2803 ), .E(\U1/aes_core/SB3/n2802 ), .F(
        \U1/aes_core/SB3/n2801 ), .Y(\U1/aes_core/SB3/n2807 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U230  ( .A(\U1/aes_core/SB3/n2807 ), .Y(
        \U1/aes_core/SB3/n2906 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U229  ( .A0(\U1/aes_core/SB3/n2875 ), 
        .A1(\U1/aes_core/SB3/n2918 ), .B0(\U1/aes_core/SB3/n2958 ), .B1(
        \U1/aes_core/SB3/n2957 ), .Y(\U1/aes_core/SB3/n2808 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U228  ( .A0(\U1/aes_core/SB3/n2865 ), 
        .A1(\U1/aes_core/SB3/n2809 ), .B0(\U1/aes_core/SB3/n2910 ), .B1(
        \U1/aes_core/SB3/n2932 ), .C0(\U1/aes_core/SB3/n2808 ), .Y(
        \U1/aes_core/SB3/n2810 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U227  ( .AN(\U1/aes_core/SB3/n2812 ), 
        .B(\U1/aes_core/SB3/n2811 ), .C(\U1/aes_core/SB3/n2906 ), .D(
        \U1/aes_core/SB3/n2810 ), .Y(\U1/aes_core/SB3/n2813 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U226  ( .A(\U1/aes_core/SB3/n2818 ), .B(
        \U1/aes_core/SB3/n2817 ), .C(\U1/aes_core/SB3/n2816 ), .D(
        \U1/aes_core/SB3/n2815 ), .E(\U1/aes_core/SB3/n2814 ), .F(
        \U1/aes_core/SB3/n2813 ), .Y(\U1/aes_core/SB3/n2883 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U225  ( .A(\U1/aes_core/SB3/n2819 ), .Y(
        \U1/aes_core/SB3/n2823 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U224  ( .A0(\U1/aes_core/SB3/n2821 ), 
        .A1(\U1/aes_core/SB3/n2820 ), .B0(\U1/aes_core/SB3/n2867 ), .B1(
        \U1/aes_core/SB3/n2826 ), .Y(\U1/aes_core/SB3/n2822 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U223  ( .A0(\U1/aes_core/SB3/n2937 ), 
        .A1(\U1/aes_core/SB3/n2824 ), .B0(\U1/aes_core/SB3/n2823 ), .C0(
        \U1/aes_core/SB3/n2822 ), .Y(\U1/aes_core/SB3/n2838 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U222  ( .A0(\U1/aes_core/SB3/n2825 ), 
        .A1(\U1/aes_core/SB3/n2909 ), .B0(\U1/aes_core/SB3/n2938 ), .Y(
        \U1/aes_core/SB3/n2830 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U221  ( .A0(\U1/aes_core/SB3/n2826 ), 
        .A1(\U1/aes_core/SB3/n2912 ), .B0(\U1/aes_core/SB3/n2941 ), .Y(
        \U1/aes_core/SB3/n2829 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U220  ( .A(\U1/aes_core/SB3/n2830 ), .B(
        \U1/aes_core/SB3/n2829 ), .C(\U1/aes_core/SB3/n2828 ), .D(
        \U1/aes_core/SB3/n2827 ), .Y(\U1/aes_core/SB3/n2837 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U219  ( .A(\U1/aes_core/SB3/n2868 ), .B(
        \U1/aes_core/SB3/n2831 ), .Y(\U1/aes_core/SB3/n2835 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U218  ( .A(\U1/aes_core/SB3/n2832 ), .B(
        \U1/aes_core/SB3/n2873 ), .Y(\U1/aes_core/SB3/n2834 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U217  ( .A0(\U1/aes_core/SB3/n2835 ), 
        .A1(\U1/aes_core/SB3/n2955 ), .B0(\U1/aes_core/SB3/n2834 ), .B1(
        \U1/aes_core/SB3/n2919 ), .C0(\U1/aes_core/SB3/n2833 ), .C1(
        \U1/aes_core/SB3/n2920 ), .Y(\U1/aes_core/SB3/n2836 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U216  ( .A(\U1/aes_core/SB3/n2928 ), .B(
        \U1/aes_core/SB3/n2883 ), .C(\U1/aes_core/SB3/n2839 ), .D(
        \U1/aes_core/SB3/n2838 ), .E(\U1/aes_core/SB3/n2837 ), .F(
        \U1/aes_core/SB3/n2836 ), .Y(\U1/aes_core/sb3 [28]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U215  ( .A1N(\U1/aes_core/SB3/n2841 ), 
        .A0(\U1/aes_core/SB3/n2840 ), .B0(\U1/aes_core/SB3/n2918 ), .Y(
        \U1/aes_core/SB3/n2857 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U214  ( .A(\U1/aes_core/SB3/n2931 ), .B(
        \U1/aes_core/SB3/n2912 ), .Y(\U1/aes_core/SB3/n2844 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U213  ( .A0(\U1/aes_core/SB3/n2955 ), 
        .A1(\U1/aes_core/SB3/n2845 ), .B0(\U1/aes_core/SB3/n2844 ), .B1(
        \U1/aes_core/SB3/n2958 ), .C0(\U1/aes_core/SB3/n2843 ), .C1(
        \U1/aes_core/SB3/n2842 ), .Y(\U1/aes_core/SB3/n2856 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U212  ( .A(\U1/aes_core/SB3/n2846 ), .Y(
        \U1/aes_core/SB3/n2849 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U211  ( .AN(\U1/aes_core/SB3/n2850 ), 
        .B(\U1/aes_core/SB3/n2849 ), .C(\U1/aes_core/SB3/n2848 ), .D(
        \U1/aes_core/SB3/n2847 ), .Y(\U1/aes_core/SB3/n2855 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U210  ( .A(\U1/aes_core/SB3/n2853 ), .B(
        \U1/aes_core/SB3/n2852 ), .C(\U1/aes_core/SB3/n2851 ), .Y(
        \U1/aes_core/SB3/n2854 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U209  ( .A(\U1/aes_core/SB3/n2859 ), .B(
        \U1/aes_core/SB3/n2858 ), .C(\U1/aes_core/SB3/n2857 ), .D(
        \U1/aes_core/SB3/n2856 ), .E(\U1/aes_core/SB3/n2855 ), .F(
        \U1/aes_core/SB3/n2854 ), .Y(\U1/aes_core/SB3/n2929 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U208  ( .A(\U1/aes_core/SB3/n2860 ), .Y(
        \U1/aes_core/SB3/n2862 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U207  ( .A0(\U1/aes_core/SB3/n2942 ), 
        .A1(\U1/aes_core/SB3/n2939 ), .B0(\U1/aes_core/SB3/n2943 ), .B1(
        \U1/aes_core/SB3/n2941 ), .Y(\U1/aes_core/SB3/n2861 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U206  ( .A0(\U1/aes_core/SB3/n2918 ), 
        .A1(\U1/aes_core/SB3/n2863 ), .B0(\U1/aes_core/SB3/n2862 ), .C0(
        \U1/aes_core/SB3/n2861 ), .Y(\U1/aes_core/SB3/n2882 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U205  ( .A0(\U1/aes_core/SB3/n2865 ), 
        .A1(\U1/aes_core/SB3/n2942 ), .B0(\U1/aes_core/SB3/n2864 ), .Y(
        \U1/aes_core/SB3/n2871 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U204  ( .A0(\U1/aes_core/SB3/n2868 ), 
        .A1(\U1/aes_core/SB3/n2867 ), .B0(\U1/aes_core/SB3/n2866 ), .Y(
        \U1/aes_core/SB3/n2870 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U203  ( .AN(\U1/aes_core/SB3/n2872 ), 
        .B(\U1/aes_core/SB3/n2871 ), .C(\U1/aes_core/SB3/n2870 ), .D(
        \U1/aes_core/SB3/n2869 ), .Y(\U1/aes_core/SB3/n2881 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U202  ( .A0(\U1/aes_core/SB3/n2938 ), 
        .A1(\U1/aes_core/SB3/n2874 ), .B0(\U1/aes_core/SB3/n2873 ), .Y(
        \U1/aes_core/SB3/n2878 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB3/U201  ( .A0(\U1/aes_core/SB3/n2920 ), .A1(
        \U1/aes_core/SB3/n2876 ), .B0(\U1/aes_core/SB3/n2957 ), .B1(
        \U1/aes_core/SB3/n2875 ), .Y(\U1/aes_core/SB3/n2877 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U200  ( .A0(\U1/aes_core/SB3/n2879 ), 
        .A1(\U1/aes_core/SB3/n2919 ), .B0(\U1/aes_core/SB3/n2878 ), .C0(
        \U1/aes_core/SB3/n2877 ), .Y(\U1/aes_core/SB3/n2880 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U199  ( .A(\U1/aes_core/SB3/n2929 ), .B(
        \U1/aes_core/SB3/n2884 ), .C(\U1/aes_core/SB3/n2883 ), .D(
        \U1/aes_core/SB3/n2882 ), .E(\U1/aes_core/SB3/n2881 ), .F(
        \U1/aes_core/SB3/n2880 ), .Y(\U1/aes_core/sb3 [29]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U198  ( .A0(\U1/aes_core/SB3/n3212 ), 
        .A1(\U1/aes_core/SB3/n3232 ), .B0(\U1/aes_core/SB3/n3253 ), .B1(
        \U1/aes_core/SB3/n3243 ), .Y(\U1/aes_core/SB3/n2885 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U197  ( .A0(\U1/aes_core/SB3/n3163 ), 
        .A1(\U1/aes_core/SB3/n3257 ), .B0(\U1/aes_core/SB3/n3113 ), .B1(
        \U1/aes_core/SB3/n3184 ), .C0(\U1/aes_core/SB3/n2885 ), .Y(
        \U1/aes_core/SB3/n2891 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U196  ( .A(\U1/aes_core/SB3/n3238 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3047 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U195  ( .A(\U1/aes_core/SB3/n3212 ), .B(
        \U1/aes_core/SB3/n3188 ), .Y(\U1/aes_core/SB3/n3028 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U194  ( .A(\U1/aes_core/SB3/n3232 ), .B(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n2996 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U193  ( .A(\U1/aes_core/SB3/n3152 ), .B(
        \U1/aes_core/SB3/n3195 ), .Y(\U1/aes_core/SB3/n3015 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U192  ( .A(\U1/aes_core/SB3/n3047 ), .B(
        \U1/aes_core/SB3/n3028 ), .C(\U1/aes_core/SB3/n2996 ), .D(
        \U1/aes_core/SB3/n3015 ), .Y(\U1/aes_core/SB3/n2890 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U191  ( .A(\U1/aes_core/SB3/n3258 ), .B(
        \U1/aes_core/SB3/n3236 ), .Y(\U1/aes_core/SB3/n3141 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U190  ( .A0(\U1/aes_core/SB3/n3189 ), 
        .A1(\U1/aes_core/SB3/n3141 ), .B0(\U1/aes_core/SB3/n3242 ), .Y(
        \U1/aes_core/SB3/n2888 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U189  ( .A0(\U1/aes_core/SB3/n3239 ), 
        .A1(\U1/aes_core/SB3/n3130 ), .B0(\U1/aes_core/SB3/n3142 ), .Y(
        \U1/aes_core/SB3/n2887 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U188  ( .A0(\U1/aes_core/SB3/n3147 ), 
        .A1(\U1/aes_core/SB3/n3187 ), .B0(\U1/aes_core/SB3/n3241 ), .Y(
        \U1/aes_core/SB3/n2886 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U187  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3239 ), .Y(\U1/aes_core/SB3/n3114 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U186  ( .A(\U1/aes_core/SB3/n2888 ), .B(
        \U1/aes_core/SB3/n2887 ), .C(\U1/aes_core/SB3/n2886 ), .D(
        \U1/aes_core/SB3/n3114 ), .Y(\U1/aes_core/SB3/n2889 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U185  ( .A(\U1/aes_core/SB3/n2894 ), .B(
        \U1/aes_core/SB3/n2893 ), .C(\U1/aes_core/SB3/n2892 ), .D(
        \U1/aes_core/SB3/n2891 ), .E(\U1/aes_core/SB3/n2890 ), .F(
        \U1/aes_core/SB3/n2889 ), .Y(\U1/aes_core/SB3/n3262 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U184  ( .A0(\U1/aes_core/SB3/n3068 ), 
        .A1(\U1/aes_core/SB3/n3243 ), .B0(\U1/aes_core/SB3/n3251 ), .B1(
        \U1/aes_core/SB3/n3186 ), .C0(\U1/aes_core/SB3/n3262 ), .Y(
        \U1/aes_core/SB3/n2895 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U183  ( .A(\U1/aes_core/SB3/n2895 ), .Y(
        \U1/aes_core/SB3/n2902 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U182  ( .A(\U1/aes_core/SB3/n3195 ), .B(
        \U1/aes_core/SB3/n2982 ), .Y(\U1/aes_core/SB3/n3104 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U181  ( .A1N(\U1/aes_core/SB3/n3104 ), 
        .A0(\U1/aes_core/SB3/n3213 ), .B0(\U1/aes_core/SB3/n3185 ), .Y(
        \U1/aes_core/SB3/n2898 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U180  ( .A0(\U1/aes_core/SB3/n3153 ), 
        .A1(\U1/aes_core/SB3/n3061 ), .B0(\U1/aes_core/SB3/n3212 ), .Y(
        \U1/aes_core/SB3/n2897 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U179  ( .A0(\U1/aes_core/SB3/n3239 ), 
        .A1(\U1/aes_core/SB3/n3194 ), .B0(\U1/aes_core/SB3/n3233 ), .Y(
        \U1/aes_core/SB3/n2896 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U178  ( .A(\U1/aes_core/SB3/n3210 ), .B(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n3011 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U177  ( .A(\U1/aes_core/SB3/n2898 ), .B(
        \U1/aes_core/SB3/n2897 ), .C(\U1/aes_core/SB3/n2896 ), .D(
        \U1/aes_core/SB3/n3011 ), .Y(\U1/aes_core/SB3/n2901 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U176  ( .A(\U1/aes_core/SB3/n3209 ), .B(
        \U1/aes_core/SB3/n3241 ), .Y(\U1/aes_core/SB3/n3240 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U175  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3187 ), .Y(\U1/aes_core/SB3/n2899 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U174  ( .A0(\U1/aes_core/SB3/n3240 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n2899 ), .B1(
        \U1/aes_core/SB3/n3221 ), .C0(\U1/aes_core/SB3/n3164 ), .C1(
        \U1/aes_core/SB3/n3166 ), .Y(\U1/aes_core/SB3/n2900 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U173  ( .A(\U1/aes_core/SB3/n2905 ), .B(
        \U1/aes_core/SB3/n2904 ), .C(\U1/aes_core/SB3/n2903 ), .D(
        \U1/aes_core/SB3/n2902 ), .E(\U1/aes_core/SB3/n2901 ), .F(
        \U1/aes_core/SB3/n2900 ), .Y(\U1/aes_core/sb3 [2]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U172  ( .A0(\U1/aes_core/SB3/n2908 ), 
        .A1(\U1/aes_core/SB3/n2948 ), .B0(\U1/aes_core/SB3/n2907 ), .B1(
        \U1/aes_core/SB3/n2955 ), .C0(\U1/aes_core/SB3/n2906 ), .Y(
        \U1/aes_core/SB3/n2926 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U171  ( .A0(\U1/aes_core/SB3/n2909 ), 
        .A1(\U1/aes_core/SB3/n2953 ), .B0(\U1/aes_core/SB3/n2942 ), .Y(
        \U1/aes_core/SB3/n2917 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U170  ( .A0(\U1/aes_core/SB3/n2933 ), 
        .A1(\U1/aes_core/SB3/n2910 ), .B0(\U1/aes_core/SB3/n2941 ), .Y(
        \U1/aes_core/SB3/n2916 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U169  ( .A0(\U1/aes_core/SB3/n2913 ), 
        .A1(\U1/aes_core/SB3/n2912 ), .B0(\U1/aes_core/SB3/n2911 ), .Y(
        \U1/aes_core/SB3/n2915 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U168  ( .A(\U1/aes_core/SB3/n2917 ), .B(
        \U1/aes_core/SB3/n2916 ), .C(\U1/aes_core/SB3/n2915 ), .D(
        \U1/aes_core/SB3/n2914 ), .Y(\U1/aes_core/SB3/n2925 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U167  ( .A(\U1/aes_core/SB3/n2948 ), .B(
        \U1/aes_core/SB3/n2918 ), .Y(\U1/aes_core/SB3/n2950 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U166  ( .A(\U1/aes_core/SB3/n2938 ), .B(
        \U1/aes_core/SB3/n2950 ), .Y(\U1/aes_core/SB3/n2922 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U165  ( .A0(\U1/aes_core/SB3/n2936 ), 
        .A1(\U1/aes_core/SB3/n2923 ), .B0(\U1/aes_core/SB3/n2922 ), .B1(
        \U1/aes_core/SB3/n2921 ), .C0(\U1/aes_core/SB3/n2920 ), .C1(
        \U1/aes_core/SB3/n2919 ), .Y(\U1/aes_core/SB3/n2924 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U164  ( .A(\U1/aes_core/SB3/n2929 ), .B(
        \U1/aes_core/SB3/n2928 ), .C(\U1/aes_core/SB3/n2927 ), .D(
        \U1/aes_core/SB3/n2926 ), .E(\U1/aes_core/SB3/n2925 ), .F(
        \U1/aes_core/SB3/n2924 ), .Y(\U1/aes_core/sb3 [30]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U163  ( .A0(\U1/aes_core/SB3/n2933 ), 
        .A1(\U1/aes_core/SB3/n2932 ), .B0(\U1/aes_core/SB3/n2931 ), .B1(
        \U1/aes_core/SB3/n2930 ), .Y(\U1/aes_core/SB3/n2934 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U162  ( .A0(\U1/aes_core/SB3/n2937 ), 
        .A1(\U1/aes_core/SB3/n2936 ), .B0(\U1/aes_core/SB3/n2935 ), .C0(
        \U1/aes_core/SB3/n2934 ), .Y(\U1/aes_core/SB3/n2961 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U161  ( .A1N(\U1/aes_core/SB3/n2940 ), 
        .A0(\U1/aes_core/SB3/n2939 ), .B0(\U1/aes_core/SB3/n2938 ), .Y(
        \U1/aes_core/SB3/n2947 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U160  ( .A0(\U1/aes_core/SB3/n2943 ), 
        .A1(\U1/aes_core/SB3/n2942 ), .B0(\U1/aes_core/SB3/n2941 ), .Y(
        \U1/aes_core/SB3/n2946 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U159  ( .A(\U1/aes_core/SB3/n2947 ), .B(
        \U1/aes_core/SB3/n2946 ), .C(\U1/aes_core/SB3/n2945 ), .D(
        \U1/aes_core/SB3/n2944 ), .Y(\U1/aes_core/SB3/n2960 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U158  ( .A(\U1/aes_core/SB3/n2949 ), .B(
        \U1/aes_core/SB3/n2948 ), .Y(\U1/aes_core/SB3/n2952 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U157  ( .A0(\U1/aes_core/SB3/n2953 ), 
        .A1(\U1/aes_core/SB3/n2952 ), .B0(\U1/aes_core/SB3/n2951 ), .B1(
        \U1/aes_core/SB3/n2950 ), .Y(\U1/aes_core/SB3/n2954 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U156  ( .A0(\U1/aes_core/SB3/n2958 ), 
        .A1(\U1/aes_core/SB3/n2957 ), .B0(\U1/aes_core/SB3/n2956 ), .B1(
        \U1/aes_core/SB3/n2955 ), .C0(\U1/aes_core/SB3/n2954 ), .Y(
        \U1/aes_core/SB3/n2959 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U155  ( .A(\U1/aes_core/SB3/n2964 ), .B(
        \U1/aes_core/SB3/n2963 ), .C(\U1/aes_core/SB3/n2962 ), .D(
        \U1/aes_core/SB3/n2961 ), .E(\U1/aes_core/SB3/n2960 ), .F(
        \U1/aes_core/SB3/n2959 ), .Y(\U1/aes_core/sb3 [31]) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U154  ( .A(\U1/aes_core/SB3/n3068 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3245 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U153  ( .AN(\U1/aes_core/SB3/n2967 ), 
        .B(\U1/aes_core/SB3/n2966 ), .C(\U1/aes_core/SB3/n2965 ), .D(
        \U1/aes_core/SB3/n3245 ), .Y(\U1/aes_core/SB3/n2974 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U152  ( .A0(\U1/aes_core/SB3/n2968 ), 
        .A1(\U1/aes_core/SB3/n3212 ), .B0(\U1/aes_core/SB3/n3130 ), .Y(
        \U1/aes_core/SB3/n2970 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U149  ( .A(\U1/aes_core/SB3/n3186 ), .B(
        \U1/aes_core/SB3/n3233 ), .Y(\U1/aes_core/SB3/n3197 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U148  ( .A0(\U1/aes_core/SB3/n3076 ), 
        .A1(\U1/aes_core/SB3/n3255 ), .B0(\U1/aes_core/SB3/n3197 ), .B1(
        \U1/aes_core/SB3/n3208 ), .C0(\U1/aes_core/SB3/n3249 ), .C1(
        \U1/aes_core/SB3/n3258 ), .Y(\U1/aes_core/SB3/n2972 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U147  ( .A(\U1/aes_core/SB3/n2977 ), .B(
        \U1/aes_core/SB3/n2976 ), .C(\U1/aes_core/SB3/n2975 ), .D(
        \U1/aes_core/SB3/n2974 ), .E(\U1/aes_core/SB3/n2973 ), .F(
        \U1/aes_core/SB3/n2972 ), .Y(\U1/aes_core/SB3/n3160 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U146  ( .AN(\U1/aes_core/SB3/n2981 ), 
        .B(\U1/aes_core/SB3/n2980 ), .C(\U1/aes_core/SB3/n2979 ), .D(
        \U1/aes_core/SB3/n2978 ), .Y(\U1/aes_core/SB3/n2991 ) );
  AOI222_X0P5M_A12TL \U1/aes_core/SB3/U145  ( .A0(\U1/aes_core/SB3/n3243 ), 
        .A1(\U1/aes_core/SB3/n3153 ), .B0(\U1/aes_core/SB3/n3238 ), .B1(
        \U1/aes_core/SB3/n3152 ), .C0(\U1/aes_core/SB3/n2982 ), .C1(
        \U1/aes_core/SB3/n3253 ), .Y(\U1/aes_core/SB3/n2990 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U144  ( .A0(\U1/aes_core/SB3/n3207 ), 
        .A1(\U1/aes_core/SB3/n3113 ), .B0(\U1/aes_core/SB3/n2983 ), .B1(
        \U1/aes_core/SB3/n3076 ), .Y(\U1/aes_core/SB3/n2984 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U143  ( .A0(\U1/aes_core/SB3/n3130 ), 
        .A1(\U1/aes_core/SB3/n3147 ), .B0(\U1/aes_core/SB3/n3146 ), .B1(
        \U1/aes_core/SB3/n3210 ), .C0(\U1/aes_core/SB3/n2984 ), .Y(
        \U1/aes_core/SB3/n2989 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U142  ( .A(\U1/aes_core/SB3/n3218 ), .B(
        \U1/aes_core/SB3/n3257 ), .Y(\U1/aes_core/SB3/n2986 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U141  ( .A0(\U1/aes_core/SB3/n3068 ), 
        .A1(\U1/aes_core/SB3/n2987 ), .B0(\U1/aes_core/SB3/n3239 ), .B1(
        \U1/aes_core/SB3/n2986 ), .C0(\U1/aes_core/SB3/n2985 ), .Y(
        \U1/aes_core/SB3/n2988 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U140  ( .AN(\U1/aes_core/SB3/n2991 ), 
        .B(\U1/aes_core/SB3/n2990 ), .C(\U1/aes_core/SB3/n2989 ), .D(
        \U1/aes_core/SB3/n2988 ), .Y(\U1/aes_core/SB3/n3205 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U139  ( .A(\U1/aes_core/SB3/n2992 ), .Y(
        \U1/aes_core/SB3/n3008 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U138  ( .A0(\U1/aes_core/SB3/n3097 ), 
        .A1(\U1/aes_core/SB3/n3166 ), .B0(\U1/aes_core/SB3/n2993 ), .Y(
        \U1/aes_core/SB3/n3007 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U137  ( .A0(\U1/aes_core/SB3/n3239 ), 
        .A1(\U1/aes_core/SB3/n3238 ), .B0(\U1/aes_core/SB3/n3209 ), .B1(
        \U1/aes_core/SB3/n2994 ), .Y(\U1/aes_core/SB3/n2995 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U136  ( .A0(\U1/aes_core/SB3/n3220 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3236 ), .B1(
        \U1/aes_core/SB3/n3248 ), .C0(\U1/aes_core/SB3/n2995 ), .Y(
        \U1/aes_core/SB3/n3006 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U135  ( .A(\U1/aes_core/SB3/n2999 ), .B(
        \U1/aes_core/SB3/n2998 ), .C(\U1/aes_core/SB3/n2997 ), .D(
        \U1/aes_core/SB3/n2996 ), .Y(\U1/aes_core/SB3/n3005 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U134  ( .AN(\U1/aes_core/SB3/n3003 ), 
        .B(\U1/aes_core/SB3/n3002 ), .C(\U1/aes_core/SB3/n3001 ), .D(
        \U1/aes_core/SB3/n3000 ), .Y(\U1/aes_core/SB3/n3004 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U133  ( .A(\U1/aes_core/SB3/n3009 ), .B(
        \U1/aes_core/SB3/n3008 ), .C(\U1/aes_core/SB3/n3007 ), .D(
        \U1/aes_core/SB3/n3006 ), .E(\U1/aes_core/SB3/n3005 ), .F(
        \U1/aes_core/SB3/n3004 ), .Y(\U1/aes_core/SB3/n3109 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U132  ( .A0(\U1/aes_core/SB3/n3196 ), 
        .A1(\U1/aes_core/SB3/n3113 ), .B0(\U1/aes_core/SB3/n3010 ), .Y(
        \U1/aes_core/SB3/n3025 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U131  ( .AN(\U1/aes_core/SB3/n3014 ), 
        .B(\U1/aes_core/SB3/n3013 ), .C(\U1/aes_core/SB3/n3012 ), .D(
        \U1/aes_core/SB3/n3011 ), .Y(\U1/aes_core/SB3/n3024 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U130  ( .A(\U1/aes_core/SB3/n3230 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3244 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U129  ( .A(\U1/aes_core/SB3/n3017 ), .B(
        \U1/aes_core/SB3/n3016 ), .C(\U1/aes_core/SB3/n3015 ), .D(
        \U1/aes_core/SB3/n3244 ), .Y(\U1/aes_core/SB3/n3023 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U128  ( .A(\U1/aes_core/SB3/n3021 ), .B(
        \U1/aes_core/SB3/n3020 ), .C(\U1/aes_core/SB3/n3019 ), .D(
        \U1/aes_core/SB3/n3018 ), .Y(\U1/aes_core/SB3/n3022 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U127  ( .A(\U1/aes_core/SB3/n3027 ), .B(
        \U1/aes_core/SB3/n3026 ), .C(\U1/aes_core/SB3/n3025 ), .D(
        \U1/aes_core/SB3/n3024 ), .E(\U1/aes_core/SB3/n3023 ), .F(
        \U1/aes_core/SB3/n3022 ), .Y(\U1/aes_core/SB3/n3133 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U126  ( .AN(\U1/aes_core/SB3/n3031 ), 
        .B(\U1/aes_core/SB3/n3030 ), .C(\U1/aes_core/SB3/n3029 ), .D(
        \U1/aes_core/SB3/n3028 ), .Y(\U1/aes_core/SB3/n3040 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U125  ( .A(\U1/aes_core/SB3/n3035 ), .B(
        \U1/aes_core/SB3/n3034 ), .C(\U1/aes_core/SB3/n3033 ), .D(
        \U1/aes_core/SB3/n3032 ), .Y(\U1/aes_core/SB3/n3039 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U124  ( .A(\U1/aes_core/SB3/n3195 ), .B(
        \U1/aes_core/SB3/n3231 ), .C(\U1/aes_core/SB3/n3233 ), .Y(
        \U1/aes_core/SB3/n3037 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U123  ( .A0(\U1/aes_core/SB3/n3037 ), 
        .A1(\U1/aes_core/SB3/n3221 ), .B0(\U1/aes_core/SB3/n3076 ), .B1(
        \U1/aes_core/SB3/n3257 ), .C0(\U1/aes_core/SB3/n3036 ), .Y(
        \U1/aes_core/SB3/n3038 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U122  ( .A(\U1/aes_core/SB3/n3043 ), .B(
        \U1/aes_core/SB3/n3042 ), .C(\U1/aes_core/SB3/n3041 ), .D(
        \U1/aes_core/SB3/n3040 ), .E(\U1/aes_core/SB3/n3039 ), .F(
        \U1/aes_core/SB3/n3038 ), .Y(\U1/aes_core/SB3/n3181 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U121  ( .A0(\U1/aes_core/SB3/n3076 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3044 ), .Y(
        \U1/aes_core/SB3/n3058 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U120  ( .A0(\U1/aes_core/SB3/n3185 ), 
        .A1(\U1/aes_core/SB3/n3187 ), .B0(\U1/aes_core/SB3/n3242 ), .B1(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3045 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U119  ( .A0(\U1/aes_core/SB3/n3096 ), 
        .A1(\U1/aes_core/SB3/n3184 ), .B0(\U1/aes_core/SB3/n3097 ), .B1(
        \U1/aes_core/SB3/n3161 ), .C0(\U1/aes_core/SB3/n3045 ), .Y(
        \U1/aes_core/SB3/n3057 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U118  ( .A(\U1/aes_core/SB3/n3046 ), .Y(
        \U1/aes_core/SB3/n3049 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U117  ( .AN(\U1/aes_core/SB3/n3050 ), 
        .B(\U1/aes_core/SB3/n3049 ), .C(\U1/aes_core/SB3/n3048 ), .D(
        \U1/aes_core/SB3/n3047 ), .Y(\U1/aes_core/SB3/n3056 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U116  ( .A(\U1/aes_core/SB3/n3054 ), .B(
        \U1/aes_core/SB3/n3053 ), .C(\U1/aes_core/SB3/n3052 ), .D(
        \U1/aes_core/SB3/n3051 ), .Y(\U1/aes_core/SB3/n3055 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U115  ( .A(\U1/aes_core/SB3/n3060 ), .B(
        \U1/aes_core/SB3/n3059 ), .C(\U1/aes_core/SB3/n3058 ), .D(
        \U1/aes_core/SB3/n3057 ), .E(\U1/aes_core/SB3/n3056 ), .F(
        \U1/aes_core/SB3/n3055 ), .Y(\U1/aes_core/SB3/n3140 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U114  ( .A0(\U1/aes_core/SB3/n3231 ), 
        .A1(\U1/aes_core/SB3/n3061 ), .B0(\U1/aes_core/SB3/n3241 ), .B1(
        \U1/aes_core/SB3/n3187 ), .Y(\U1/aes_core/SB3/n3062 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U113  ( .A0(\U1/aes_core/SB3/n3113 ), 
        .A1(\U1/aes_core/SB3/n3258 ), .B0(\U1/aes_core/SB3/n3063 ), .B1(
        \U1/aes_core/SB3/n3248 ), .C0(\U1/aes_core/SB3/n3062 ), .Y(
        \U1/aes_core/SB3/n3075 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U112  ( .AN(\U1/aes_core/SB3/n3067 ), 
        .B(\U1/aes_core/SB3/n3066 ), .C(\U1/aes_core/SB3/n3065 ), .D(
        \U1/aes_core/SB3/n3064 ), .Y(\U1/aes_core/SB3/n3074 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U111  ( .A0(\U1/aes_core/SB3/n3251 ), 
        .A1(\U1/aes_core/SB3/n3068 ), .B0(\U1/aes_core/SB3/n3242 ), .Y(
        \U1/aes_core/SB3/n3072 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U110  ( .A(\U1/aes_core/SB3/n3218 ), .B(
        \U1/aes_core/SB3/n3223 ), .Y(\U1/aes_core/SB3/n3069 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U109  ( .A0(\U1/aes_core/SB3/n3194 ), 
        .A1(\U1/aes_core/SB3/n3069 ), .B0(\U1/aes_core/SB3/n3195 ), .B1(
        \U1/aes_core/SB3/n3141 ), .Y(\U1/aes_core/SB3/n3070 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U108  ( .A(\U1/aes_core/SB3/n3072 ), .B(
        \U1/aes_core/SB3/n3071 ), .C(\U1/aes_core/SB3/n3070 ), .Y(
        \U1/aes_core/SB3/n3073 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U107  ( .A(\U1/aes_core/SB3/n3133 ), .B(
        \U1/aes_core/SB3/n3181 ), .C(\U1/aes_core/SB3/n3140 ), .D(
        \U1/aes_core/SB3/n3075 ), .E(\U1/aes_core/SB3/n3074 ), .F(
        \U1/aes_core/SB3/n3073 ), .Y(\U1/aes_core/SB3/n3227 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U106  ( .A(\U1/aes_core/SB3/n3160 ), .B(
        \U1/aes_core/SB3/n3205 ), .C(\U1/aes_core/SB3/n3109 ), .D(
        \U1/aes_core/SB3/n3227 ), .Y(\U1/aes_core/SB3/n3089 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U105  ( .A0(\U1/aes_core/SB3/n3207 ), 
        .A1(\U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3076 ), .B1(
        \U1/aes_core/SB3/n3223 ), .Y(\U1/aes_core/SB3/n3077 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U104  ( .A0(\U1/aes_core/SB3/n3212 ), 
        .A1(\U1/aes_core/SB3/n3230 ), .B0(\U1/aes_core/SB3/n3243 ), .B1(
        \U1/aes_core/SB3/n3251 ), .C0(\U1/aes_core/SB3/n3077 ), .Y(
        \U1/aes_core/SB3/n3088 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U103  ( .A(\U1/aes_core/SB3/n3078 ), .Y(
        \U1/aes_core/SB3/n3081 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U102  ( .A0(\U1/aes_core/SB3/n3079 ), 
        .A1(\U1/aes_core/SB3/n3184 ), .B0(\U1/aes_core/SB3/n3112 ), .B1(
        \U1/aes_core/SB3/n3164 ), .Y(\U1/aes_core/SB3/n3080 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U101  ( .A0(\U1/aes_core/SB3/n3231 ), 
        .A1(\U1/aes_core/SB3/n3081 ), .B0(\U1/aes_core/SB3/n3213 ), .B1(
        \U1/aes_core/SB3/n3162 ), .C0(\U1/aes_core/SB3/n3080 ), .Y(
        \U1/aes_core/SB3/n3087 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U100  ( .A0(\U1/aes_core/SB3/n3253 ), 
        .A1(\U1/aes_core/SB3/n3130 ), .B0(\U1/aes_core/SB3/n3233 ), .Y(
        \U1/aes_core/SB3/n3085 ) );
  AND4_X0P5M_A12TL \U1/aes_core/SB3/U99  ( .A(\U1/aes_core/SB3/n3085 ), .B(
        \U1/aes_core/SB3/n3084 ), .C(\U1/aes_core/SB3/n3083 ), .D(
        \U1/aes_core/SB3/n3082 ), .Y(\U1/aes_core/SB3/n3086 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U98  ( .AN(\U1/aes_core/SB3/n3089 ), .B(
        \U1/aes_core/SB3/n3088 ), .C(\U1/aes_core/SB3/n3087 ), .D(
        \U1/aes_core/SB3/n3086 ), .Y(\U1/aes_core/sb3 [3]) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U97  ( .A0(\U1/aes_core/SB3/n3104 ), .A1(
        \U1/aes_core/SB3/n3219 ), .B0(\U1/aes_core/SB3/n3163 ), .Y(
        \U1/aes_core/SB3/n3101 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U96  ( .A(\U1/aes_core/SB3/n3092 ), .B(
        \U1/aes_core/SB3/n3091 ), .C(\U1/aes_core/SB3/n3090 ), .Y(
        \U1/aes_core/SB3/n3100 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U95  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3242 ), .Y(\U1/aes_core/SB3/n3095 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U94  ( .A(\U1/aes_core/SB3/n3213 ), .B(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3093 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U93  ( .A0(\U1/aes_core/SB3/n3095 ), 
        .A1(\U1/aes_core/SB3/n3094 ), .B0(\U1/aes_core/SB3/n3093 ), .B1(
        \U1/aes_core/SB3/n3236 ), .C0(\U1/aes_core/SB3/n3219 ), .C1(
        \U1/aes_core/SB3/n3145 ), .Y(\U1/aes_core/SB3/n3099 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U92  ( .A0(\U1/aes_core/SB3/n3196 ), 
        .A1(\U1/aes_core/SB3/n3097 ), .B0(\U1/aes_core/SB3/n3258 ), .B1(
        \U1/aes_core/SB3/n3248 ), .C0(\U1/aes_core/SB3/n3221 ), .C1(
        \U1/aes_core/SB3/n3096 ), .Y(\U1/aes_core/SB3/n3098 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U91  ( .A(\U1/aes_core/SB3/n3103 ), .B(
        \U1/aes_core/SB3/n3102 ), .C(\U1/aes_core/SB3/n3101 ), .D(
        \U1/aes_core/SB3/n3100 ), .E(\U1/aes_core/SB3/n3099 ), .F(
        \U1/aes_core/SB3/n3098 ), .Y(\U1/aes_core/SB3/n3228 ) );
  AOI21_X0P5M_A12TL \U1/aes_core/SB3/U90  ( .A0(\U1/aes_core/SB3/n3104 ), .A1(
        \U1/aes_core/SB3/n3113 ), .B0(\U1/aes_core/SB3/n3184 ), .Y(
        \U1/aes_core/SB3/n3139 ) );
  AOI31_X0P5M_A12TL \U1/aes_core/SB3/U89  ( .A0(\U1/aes_core/SB3/n3208 ), .A1(
        \U1/aes_core/SB3/n3221 ), .A2(\U1/aes_core/SB3/n3161 ), .B0(
        \U1/aes_core/SB3/n3237 ), .Y(\U1/aes_core/SB3/n3138 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U88  ( .A(\U1/aes_core/SB3/n3108 ), .B(
        \U1/aes_core/SB3/n3107 ), .C(\U1/aes_core/SB3/n3106 ), .D(
        \U1/aes_core/SB3/n3105 ), .Y(\U1/aes_core/SB3/n3135 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U87  ( .A(\U1/aes_core/SB3/n3109 ), .Y(
        \U1/aes_core/SB3/n3132 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U86  ( .A(\U1/aes_core/SB3/n3110 ), .Y(
        \U1/aes_core/SB3/n3126 ) );
  OAI21B_X0P5M_A12TL \U1/aes_core/SB3/U85  ( .A0(\U1/aes_core/SB3/n3112 ), 
        .A1(\U1/aes_core/SB3/n3249 ), .B0N(\U1/aes_core/SB3/n3111 ), .Y(
        \U1/aes_core/SB3/n3125 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U84  ( .A0(\U1/aes_core/SB3/n3256 ), 
        .A1(\U1/aes_core/SB3/n3113 ), .B0(\U1/aes_core/SB3/n3163 ), .B1(
        \U1/aes_core/SB3/n3223 ), .C0(\U1/aes_core/SB3/n3237 ), .C1(
        \U1/aes_core/SB3/n3258 ), .Y(\U1/aes_core/SB3/n3124 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U83  ( .AN(\U1/aes_core/SB3/n3117 ), .B(
        \U1/aes_core/SB3/n3116 ), .C(\U1/aes_core/SB3/n3115 ), .D(
        \U1/aes_core/SB3/n3114 ), .Y(\U1/aes_core/SB3/n3123 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U82  ( .A(\U1/aes_core/SB3/n3121 ), .B(
        \U1/aes_core/SB3/n3120 ), .C(\U1/aes_core/SB3/n3119 ), .D(
        \U1/aes_core/SB3/n3118 ), .Y(\U1/aes_core/SB3/n3122 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U81  ( .A(\U1/aes_core/SB3/n3127 ), .B(
        \U1/aes_core/SB3/n3126 ), .C(\U1/aes_core/SB3/n3125 ), .D(
        \U1/aes_core/SB3/n3124 ), .E(\U1/aes_core/SB3/n3123 ), .F(
        \U1/aes_core/SB3/n3122 ), .Y(\U1/aes_core/SB3/n3128 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U80  ( .A(\U1/aes_core/SB3/n3128 ), .Y(
        \U1/aes_core/SB3/n3206 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U79  ( .A0(\U1/aes_core/SB3/n3196 ), .A1(
        \U1/aes_core/SB3/n3218 ), .B0(\U1/aes_core/SB3/n3258 ), .B1(
        \U1/aes_core/SB3/n3257 ), .Y(\U1/aes_core/SB3/n3129 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U78  ( .A0(\U1/aes_core/SB3/n3186 ), 
        .A1(\U1/aes_core/SB3/n3130 ), .B0(\U1/aes_core/SB3/n3210 ), .B1(
        \U1/aes_core/SB3/n3232 ), .C0(\U1/aes_core/SB3/n3129 ), .Y(
        \U1/aes_core/SB3/n3131 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U77  ( .AN(\U1/aes_core/SB3/n3133 ), .B(
        \U1/aes_core/SB3/n3132 ), .C(\U1/aes_core/SB3/n3206 ), .D(
        \U1/aes_core/SB3/n3131 ), .Y(\U1/aes_core/SB3/n3134 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U76  ( .A(\U1/aes_core/SB3/n3139 ), .B(
        \U1/aes_core/SB3/n3138 ), .C(\U1/aes_core/SB3/n3137 ), .D(
        \U1/aes_core/SB3/n3136 ), .E(\U1/aes_core/SB3/n3135 ), .F(
        \U1/aes_core/SB3/n3134 ), .Y(\U1/aes_core/SB3/n3204 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U75  ( .A(\U1/aes_core/SB3/n3140 ), .Y(
        \U1/aes_core/SB3/n3144 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U74  ( .A0(\U1/aes_core/SB3/n3142 ), .A1(
        \U1/aes_core/SB3/n3141 ), .B0(\U1/aes_core/SB3/n3188 ), .B1(
        \U1/aes_core/SB3/n3147 ), .Y(\U1/aes_core/SB3/n3143 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U73  ( .A0(\U1/aes_core/SB3/n3237 ), 
        .A1(\U1/aes_core/SB3/n3145 ), .B0(\U1/aes_core/SB3/n3144 ), .C0(
        \U1/aes_core/SB3/n3143 ), .Y(\U1/aes_core/SB3/n3159 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U72  ( .A0(\U1/aes_core/SB3/n3146 ), .A1(
        \U1/aes_core/SB3/n3209 ), .B0(\U1/aes_core/SB3/n3238 ), .Y(
        \U1/aes_core/SB3/n3151 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U71  ( .A0(\U1/aes_core/SB3/n3147 ), .A1(
        \U1/aes_core/SB3/n3212 ), .B0(\U1/aes_core/SB3/n3241 ), .Y(
        \U1/aes_core/SB3/n3150 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U70  ( .A(\U1/aes_core/SB3/n3151 ), .B(
        \U1/aes_core/SB3/n3150 ), .C(\U1/aes_core/SB3/n3149 ), .D(
        \U1/aes_core/SB3/n3148 ), .Y(\U1/aes_core/SB3/n3158 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U69  ( .A(\U1/aes_core/SB3/n3189 ), .B(
        \U1/aes_core/SB3/n3152 ), .Y(\U1/aes_core/SB3/n3156 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U68  ( .A(\U1/aes_core/SB3/n3153 ), .B(
        \U1/aes_core/SB3/n3194 ), .Y(\U1/aes_core/SB3/n3155 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U67  ( .A0(\U1/aes_core/SB3/n3156 ), 
        .A1(\U1/aes_core/SB3/n3255 ), .B0(\U1/aes_core/SB3/n3155 ), .B1(
        \U1/aes_core/SB3/n3219 ), .C0(\U1/aes_core/SB3/n3154 ), .C1(
        \U1/aes_core/SB3/n3220 ), .Y(\U1/aes_core/SB3/n3157 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U66  ( .A(\U1/aes_core/SB3/n3228 ), .B(
        \U1/aes_core/SB3/n3204 ), .C(\U1/aes_core/SB3/n3160 ), .D(
        \U1/aes_core/SB3/n3159 ), .E(\U1/aes_core/SB3/n3158 ), .F(
        \U1/aes_core/SB3/n3157 ), .Y(\U1/aes_core/sb3 [4]) );
  AOI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U65  ( .A1N(\U1/aes_core/SB3/n3162 ), 
        .A0(\U1/aes_core/SB3/n3161 ), .B0(\U1/aes_core/SB3/n3218 ), .Y(
        \U1/aes_core/SB3/n3178 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U64  ( .A(\U1/aes_core/SB3/n3231 ), .B(
        \U1/aes_core/SB3/n3212 ), .Y(\U1/aes_core/SB3/n3165 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U63  ( .A0(\U1/aes_core/SB3/n3255 ), 
        .A1(\U1/aes_core/SB3/n3166 ), .B0(\U1/aes_core/SB3/n3165 ), .B1(
        \U1/aes_core/SB3/n3258 ), .C0(\U1/aes_core/SB3/n3164 ), .C1(
        \U1/aes_core/SB3/n3163 ), .Y(\U1/aes_core/SB3/n3177 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U62  ( .A(\U1/aes_core/SB3/n3167 ), .Y(
        \U1/aes_core/SB3/n3170 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U61  ( .AN(\U1/aes_core/SB3/n3171 ), .B(
        \U1/aes_core/SB3/n3170 ), .C(\U1/aes_core/SB3/n3169 ), .D(
        \U1/aes_core/SB3/n3168 ), .Y(\U1/aes_core/SB3/n3176 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U60  ( .A(\U1/aes_core/SB3/n3174 ), .B(
        \U1/aes_core/SB3/n3173 ), .C(\U1/aes_core/SB3/n3172 ), .Y(
        \U1/aes_core/SB3/n3175 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U59  ( .A(\U1/aes_core/SB3/n3180 ), .B(
        \U1/aes_core/SB3/n3179 ), .C(\U1/aes_core/SB3/n3178 ), .D(
        \U1/aes_core/SB3/n3177 ), .E(\U1/aes_core/SB3/n3176 ), .F(
        \U1/aes_core/SB3/n3175 ), .Y(\U1/aes_core/SB3/n3229 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U58  ( .A(\U1/aes_core/SB3/n3181 ), .Y(
        \U1/aes_core/SB3/n3183 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U57  ( .A0(\U1/aes_core/SB3/n3242 ), .A1(
        \U1/aes_core/SB3/n3239 ), .B0(\U1/aes_core/SB3/n3243 ), .B1(
        \U1/aes_core/SB3/n3241 ), .Y(\U1/aes_core/SB3/n3182 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U56  ( .A0(\U1/aes_core/SB3/n3218 ), 
        .A1(\U1/aes_core/SB3/n3184 ), .B0(\U1/aes_core/SB3/n3183 ), .C0(
        \U1/aes_core/SB3/n3182 ), .Y(\U1/aes_core/SB3/n3203 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U55  ( .A0(\U1/aes_core/SB3/n3186 ), .A1(
        \U1/aes_core/SB3/n3242 ), .B0(\U1/aes_core/SB3/n3185 ), .Y(
        \U1/aes_core/SB3/n3192 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U54  ( .A0(\U1/aes_core/SB3/n3189 ), .A1(
        \U1/aes_core/SB3/n3188 ), .B0(\U1/aes_core/SB3/n3187 ), .Y(
        \U1/aes_core/SB3/n3191 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U53  ( .AN(\U1/aes_core/SB3/n3193 ), .B(
        \U1/aes_core/SB3/n3192 ), .C(\U1/aes_core/SB3/n3191 ), .D(
        \U1/aes_core/SB3/n3190 ), .Y(\U1/aes_core/SB3/n3202 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U52  ( .A0(\U1/aes_core/SB3/n3238 ), .A1(
        \U1/aes_core/SB3/n3195 ), .B0(\U1/aes_core/SB3/n3194 ), .Y(
        \U1/aes_core/SB3/n3199 ) );
  OA22_X0P5M_A12TL \U1/aes_core/SB3/U51  ( .A0(\U1/aes_core/SB3/n3220 ), .A1(
        \U1/aes_core/SB3/n3197 ), .B0(\U1/aes_core/SB3/n3257 ), .B1(
        \U1/aes_core/SB3/n3196 ), .Y(\U1/aes_core/SB3/n3198 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U50  ( .A0(\U1/aes_core/SB3/n3200 ), 
        .A1(\U1/aes_core/SB3/n3219 ), .B0(\U1/aes_core/SB3/n3199 ), .C0(
        \U1/aes_core/SB3/n3198 ), .Y(\U1/aes_core/SB3/n3201 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U49  ( .A(\U1/aes_core/SB3/n3229 ), .B(
        \U1/aes_core/SB3/n3205 ), .C(\U1/aes_core/SB3/n3204 ), .D(
        \U1/aes_core/SB3/n3203 ), .E(\U1/aes_core/SB3/n3202 ), .F(
        \U1/aes_core/SB3/n3201 ), .Y(\U1/aes_core/sb3 [5]) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U48  ( .A0(\U1/aes_core/SB3/n3208 ), 
        .A1(\U1/aes_core/SB3/n3248 ), .B0(\U1/aes_core/SB3/n3207 ), .B1(
        \U1/aes_core/SB3/n3255 ), .C0(\U1/aes_core/SB3/n3206 ), .Y(
        \U1/aes_core/SB3/n3226 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U47  ( .A0(\U1/aes_core/SB3/n3209 ), .A1(
        \U1/aes_core/SB3/n3253 ), .B0(\U1/aes_core/SB3/n3242 ), .Y(
        \U1/aes_core/SB3/n3217 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U46  ( .A0(\U1/aes_core/SB3/n3233 ), .A1(
        \U1/aes_core/SB3/n3210 ), .B0(\U1/aes_core/SB3/n3241 ), .Y(
        \U1/aes_core/SB3/n3216 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U45  ( .A0(\U1/aes_core/SB3/n3213 ), .A1(
        \U1/aes_core/SB3/n3212 ), .B0(\U1/aes_core/SB3/n3211 ), .Y(
        \U1/aes_core/SB3/n3215 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U44  ( .A(\U1/aes_core/SB3/n3217 ), .B(
        \U1/aes_core/SB3/n3216 ), .C(\U1/aes_core/SB3/n3215 ), .D(
        \U1/aes_core/SB3/n3214 ), .Y(\U1/aes_core/SB3/n3225 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U43  ( .A(\U1/aes_core/SB3/n3248 ), .B(
        \U1/aes_core/SB3/n3218 ), .Y(\U1/aes_core/SB3/n3250 ) );
  NOR2_X0P5A_A12TL \U1/aes_core/SB3/U42  ( .A(\U1/aes_core/SB3/n3238 ), .B(
        \U1/aes_core/SB3/n3250 ), .Y(\U1/aes_core/SB3/n3222 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U41  ( .A0(\U1/aes_core/SB3/n3236 ), 
        .A1(\U1/aes_core/SB3/n3223 ), .B0(\U1/aes_core/SB3/n3222 ), .B1(
        \U1/aes_core/SB3/n3221 ), .C0(\U1/aes_core/SB3/n3220 ), .C1(
        \U1/aes_core/SB3/n3219 ), .Y(\U1/aes_core/SB3/n3224 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U40  ( .A(\U1/aes_core/SB3/n3229 ), .B(
        \U1/aes_core/SB3/n3228 ), .C(\U1/aes_core/SB3/n3227 ), .D(
        \U1/aes_core/SB3/n3226 ), .E(\U1/aes_core/SB3/n3225 ), .F(
        \U1/aes_core/SB3/n3224 ), .Y(\U1/aes_core/sb3 [6]) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U39  ( .A0(\U1/aes_core/SB3/n3233 ), .A1(
        \U1/aes_core/SB3/n3232 ), .B0(\U1/aes_core/SB3/n3231 ), .B1(
        \U1/aes_core/SB3/n3230 ), .Y(\U1/aes_core/SB3/n3234 ) );
  OAI211_X0P5M_A12TL \U1/aes_core/SB3/U38  ( .A0(\U1/aes_core/SB3/n3237 ), 
        .A1(\U1/aes_core/SB3/n3236 ), .B0(\U1/aes_core/SB3/n3235 ), .C0(
        \U1/aes_core/SB3/n3234 ), .Y(\U1/aes_core/SB3/n3261 ) );
  OAI2XB1_X0P5M_A12TL \U1/aes_core/SB3/U37  ( .A1N(\U1/aes_core/SB3/n3240 ), 
        .A0(\U1/aes_core/SB3/n3239 ), .B0(\U1/aes_core/SB3/n3238 ), .Y(
        \U1/aes_core/SB3/n3247 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U36  ( .A0(\U1/aes_core/SB3/n3243 ), .A1(
        \U1/aes_core/SB3/n3242 ), .B0(\U1/aes_core/SB3/n3241 ), .Y(
        \U1/aes_core/SB3/n3246 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U35  ( .A(\U1/aes_core/SB3/n3247 ), .B(
        \U1/aes_core/SB3/n3246 ), .C(\U1/aes_core/SB3/n3245 ), .D(
        \U1/aes_core/SB3/n3244 ), .Y(\U1/aes_core/SB3/n3260 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U34  ( .A(\U1/aes_core/SB3/n3249 ), .B(
        \U1/aes_core/SB3/n3248 ), .Y(\U1/aes_core/SB3/n3252 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U33  ( .A0(\U1/aes_core/SB3/n3253 ), .A1(
        \U1/aes_core/SB3/n3252 ), .B0(\U1/aes_core/SB3/n3251 ), .B1(
        \U1/aes_core/SB3/n3250 ), .Y(\U1/aes_core/SB3/n3254 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U32  ( .A0(\U1/aes_core/SB3/n3258 ), 
        .A1(\U1/aes_core/SB3/n3257 ), .B0(\U1/aes_core/SB3/n3256 ), .B1(
        \U1/aes_core/SB3/n3255 ), .C0(\U1/aes_core/SB3/n3254 ), .Y(
        \U1/aes_core/SB3/n3259 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U31  ( .A(\U1/aes_core/SB3/n3264 ), .B(
        \U1/aes_core/SB3/n3263 ), .C(\U1/aes_core/SB3/n3262 ), .D(
        \U1/aes_core/SB3/n3261 ), .E(\U1/aes_core/SB3/n3260 ), .F(
        \U1/aes_core/SB3/n3259 ), .Y(\U1/aes_core/sb3 [7]) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U30  ( .A(\U1/aes_core/SB3/n3267 ), .B(
        \U1/aes_core/SB3/n3266 ), .C(\U1/aes_core/SB3/n3265 ), .Y(
        \U1/aes_core/SB3/n3290 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U29  ( .A0(\U1/aes_core/SB3/n3268 ), .A1(
        \U1/aes_core/SB3/n3324 ), .B0(\U1/aes_core/SB3/n3340 ), .Y(
        \U1/aes_core/SB3/n3273 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U28  ( .A0(\U1/aes_core/SB3/n3333 ), .A1(
        \U1/aes_core/SB3/n3270 ), .B0(\U1/aes_core/SB3/n3269 ), .B1(
        \U1/aes_core/SB3/n3334 ), .Y(\U1/aes_core/SB3/n3271 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U27  ( .A(\U1/aes_core/SB3/n3273 ), .B(
        \U1/aes_core/SB3/n3272 ), .C(\U1/aes_core/SB3/n3271 ), .Y(
        \U1/aes_core/SB3/n3289 ) );
  AOI22_X0P5M_A12TL \U1/aes_core/SB3/U26  ( .A0(\U1/aes_core/SB3/n3276 ), .A1(
        \U1/aes_core/SB3/n3299 ), .B0(\U1/aes_core/SB3/n3275 ), .B1(
        \U1/aes_core/SB3/n3274 ), .Y(\U1/aes_core/SB3/n3277 ) );
  OAI221_X0P5M_A12TL \U1/aes_core/SB3/U25  ( .A0(\U1/aes_core/SB3/n3281 ), 
        .A1(\U1/aes_core/SB3/n3280 ), .B0(\U1/aes_core/SB3/n3279 ), .B1(
        \U1/aes_core/SB3/n3278 ), .C0(\U1/aes_core/SB3/n3277 ), .Y(
        \U1/aes_core/SB3/n3288 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U24  ( .A(\U1/aes_core/SB3/n3329 ), .B(
        \U1/aes_core/SB3/n3282 ), .Y(\U1/aes_core/SB3/n3283 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U23  ( .AN(\U1/aes_core/SB3/n3286 ), .B(
        \U1/aes_core/SB3/n3285 ), .C(\U1/aes_core/SB3/n3284 ), .D(
        \U1/aes_core/SB3/n3283 ), .Y(\U1/aes_core/SB3/n3287 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U22  ( .A(\U1/aes_core/SB3/n3292 ), .B(
        \U1/aes_core/SB3/n3291 ), .C(\U1/aes_core/SB3/n3290 ), .D(
        \U1/aes_core/SB3/n3289 ), .E(\U1/aes_core/SB3/n3288 ), .F(
        \U1/aes_core/SB3/n3287 ), .Y(\U1/aes_core/SB3/n3351 ) );
  OR4_X0P5M_A12TL \U1/aes_core/SB3/U21  ( .A(\U1/aes_core/SB3/n3295 ), .B(
        \U1/aes_core/SB3/n3294 ), .C(\U1/aes_core/SB3/n3293 ), .D(
        \U1/aes_core/SB3/n3351 ), .Y(\U1/aes_core/SB3/n3320 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U20  ( .A0(\U1/aes_core/SB3/n3297 ), .A1(
        \U1/aes_core/SB3/n3308 ), .B0(\U1/aes_core/SB3/n3344 ), .B1(
        \U1/aes_core/SB3/n3296 ), .Y(\U1/aes_core/SB3/n3298 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U19  ( .A0(\U1/aes_core/SB3/n3322 ), 
        .A1(\U1/aes_core/SB3/n3334 ), .B0(\U1/aes_core/SB3/n3325 ), .B1(
        \U1/aes_core/SB3/n3299 ), .C0(\U1/aes_core/SB3/n3298 ), .Y(
        \U1/aes_core/SB3/n3319 ) );
  OAI22_X0P5M_A12TL \U1/aes_core/SB3/U18  ( .A0(\U1/aes_core/SB3/n3303 ), .A1(
        \U1/aes_core/SB3/n3302 ), .B0(\U1/aes_core/SB3/n3301 ), .B1(
        \U1/aes_core/SB3/n3300 ), .Y(\U1/aes_core/SB3/n3304 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U17  ( .A0(\U1/aes_core/SB3/n3307 ), 
        .A1(\U1/aes_core/SB3/n3306 ), .B0(\U1/aes_core/SB3/n3305 ), .B1(
        \U1/aes_core/SB3/n3330 ), .C0(\U1/aes_core/SB3/n3304 ), .Y(
        \U1/aes_core/SB3/n3318 ) );
  NAND2_X0P5A_A12TL \U1/aes_core/SB3/U16  ( .A(\U1/aes_core/SB3/n3309 ), .B(
        \U1/aes_core/SB3/n3308 ), .Y(\U1/aes_core/SB3/n3316 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U15  ( .A(\U1/aes_core/SB3/n3310 ), .Y(
        \U1/aes_core/SB3/n3315 ) );
  NAND3_X0P5A_A12TL \U1/aes_core/SB3/U14  ( .A(\U1/aes_core/SB3/n3313 ), .B(
        \U1/aes_core/SB3/n3312 ), .C(\U1/aes_core/SB3/n3311 ), .Y(
        \U1/aes_core/SB3/n3314 ) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U13  ( .A0(\U1/aes_core/SB3/n3331 ), 
        .A1(\U1/aes_core/SB3/n3316 ), .B0(\U1/aes_core/SB3/n3323 ), .B1(
        \U1/aes_core/SB3/n3315 ), .C0(\U1/aes_core/SB3/n3314 ), .Y(
        \U1/aes_core/SB3/n3317 ) );
  NAND4B_X0P5M_A12TL \U1/aes_core/SB3/U12  ( .AN(\U1/aes_core/SB3/n3320 ), .B(
        \U1/aes_core/SB3/n3319 ), .C(\U1/aes_core/SB3/n3318 ), .D(
        \U1/aes_core/SB3/n3317 ), .Y(\U1/aes_core/sb3 [8]) );
  AOI221_X0P5M_A12TL \U1/aes_core/SB3/U11  ( .A0(\U1/aes_core/SB3/n3325 ), 
        .A1(\U1/aes_core/SB3/n3324 ), .B0(\U1/aes_core/SB3/n3323 ), .B1(
        \U1/aes_core/SB3/n3322 ), .C0(\U1/aes_core/SB3/n3321 ), .Y(
        \U1/aes_core/SB3/n3326 ) );
  INV_X0P5B_A12TL \U1/aes_core/SB3/U10  ( .A(\U1/aes_core/SB3/n3326 ), .Y(
        \U1/aes_core/SB3/n3350 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U9  ( .A0(\U1/aes_core/SB3/n3339 ), .A1(
        \U1/aes_core/SB3/n3328 ), .B0(\U1/aes_core/SB3/n3327 ), .Y(
        \U1/aes_core/SB3/n3338 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U8  ( .A0(\U1/aes_core/SB3/n3331 ), .A1(
        \U1/aes_core/SB3/n3330 ), .B0(\U1/aes_core/SB3/n3329 ), .Y(
        \U1/aes_core/SB3/n3337 ) );
  OAI21_X0P5M_A12TL \U1/aes_core/SB3/U7  ( .A0(\U1/aes_core/SB3/n3334 ), .A1(
        \U1/aes_core/SB3/n3333 ), .B0(\U1/aes_core/SB3/n3332 ), .Y(
        \U1/aes_core/SB3/n3336 ) );
  NAND4_X0P5A_A12TL \U1/aes_core/SB3/U6  ( .A(\U1/aes_core/SB3/n3338 ), .B(
        \U1/aes_core/SB3/n3337 ), .C(\U1/aes_core/SB3/n3336 ), .D(
        \U1/aes_core/SB3/n3335 ), .Y(\U1/aes_core/SB3/n3349 ) );
  NOR3_X0P5A_A12TL \U1/aes_core/SB3/U5  ( .A(\U1/aes_core/SB3/n3341 ), .B(
        \U1/aes_core/SB3/n3340 ), .C(\U1/aes_core/SB3/n3339 ), .Y(
        \U1/aes_core/SB3/n3345 ) );
  OAI222_X0P5M_A12TL \U1/aes_core/SB3/U4  ( .A0(\U1/aes_core/SB3/n3347 ), .A1(
        \U1/aes_core/SB3/n3346 ), .B0(\U1/aes_core/SB3/n3345 ), .B1(
        \U1/aes_core/SB3/n3344 ), .C0(\U1/aes_core/SB3/n3343 ), .C1(
        \U1/aes_core/SB3/n3342 ), .Y(\U1/aes_core/SB3/n3348 ) );
  OR6_X0P5M_A12TL \U1/aes_core/SB3/U3  ( .A(\U1/aes_core/SB3/n3353 ), .B(
        \U1/aes_core/SB3/n3352 ), .C(\U1/aes_core/SB3/n3351 ), .D(
        \U1/aes_core/SB3/n3350 ), .E(\U1/aes_core/SB3/n3349 ), .F(
        \U1/aes_core/SB3/n3348 ), .Y(\U1/aes_core/sb3 [9]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U30  ( .A(\U1/aes_core/MC0/n36 ), .B(
        \U1/aes_core/MC0/n35 ), .Y(\U1/aes_core/sc0 [28]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U3  ( .A(\U1/aes_core/MC0/n23 ), .B(
        \U1/aes_core/MC0/n38 ), .Y(\U1/aes_core/sc0 [27]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U1  ( .A(\U1/aes_core/MC0/n4 ), .B(
        \U1/aes_core/MC0/n2 ), .Y(\U1/aes_core/sc0 [9]) );
  INV_X0P5B_A12TL \U1/aes_core/MC0/U112  ( .A(\U1/aes_core/sb2 [8]), .Y(
        \U1/aes_core/MC0/n66 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U111  ( .A(\U1/aes_core/MC0/n66 ), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/MC0/n79 ) );
  INV_X0P5B_A12TL \U1/aes_core/MC0/U110  ( .A(\U1/aes_core/sb0 [31]), .Y(
        \U1/aes_core/MC0/n11 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U109  ( .A(\U1/aes_core/sb1 [16]), .B(
        \U1/aes_core/MC0/n11 ), .Y(\U1/aes_core/MC0/n46 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U108  ( .A(\U1/aes_core/sb0 [24]), .B(
        \U1/aes_core/MC0/n46 ), .Y(\U1/aes_core/MC0/n80 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U107  ( .A(\U1/aes_core/MC0/n79 ), .B(
        \U1/aes_core/MC0/n80 ), .Y(\U1/aes_core/sc0 [0]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U106  ( .A(\U1/aes_core/sb0 [26]), .B(
        \U1/aes_core/sb3 [2]), .Y(\U1/aes_core/MC0/n64 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U105  ( .A(\U1/aes_core/sb3 [1]), .B(
        \U1/aes_core/sb2 [9]), .Y(\U1/aes_core/MC0/n68 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U104  ( .A(\U1/aes_core/sb1 [18]), .B(
        \U1/aes_core/MC0/n68 ), .Y(\U1/aes_core/MC0/n78 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U103  ( .A(\U1/aes_core/MC0/n64 ), .B(
        \U1/aes_core/MC0/n78 ), .Y(\U1/aes_core/sc0 [10]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U102  ( .A(\U1/aes_core/sb1 [19]), .B(
        \U1/aes_core/sb3 [3]), .Y(\U1/aes_core/MC0/n75 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U101  ( .A(\U1/aes_core/sb0 [27]), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/MC0/n77 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U100  ( .A(\U1/aes_core/MC0/n77 ), .B(
        \U1/aes_core/sb2 [10]), .Y(\U1/aes_core/MC0/n59 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U99  ( .A(\U1/aes_core/sb3 [2]), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/MC0/n24 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U98  ( .A(\U1/aes_core/MC0/n59 ), .B(
        \U1/aes_core/MC0/n24 ), .Y(\U1/aes_core/MC0/n76 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U97  ( .A(\U1/aes_core/MC0/n75 ), .B(
        \U1/aes_core/MC0/n76 ), .Y(\U1/aes_core/sc0 [11]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U96  ( .A(\U1/aes_core/sb2 [11]), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/MC0/n54 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U95  ( .A(\U1/aes_core/sb3 [3]), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/MC0/n74 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U94  ( .A(\U1/aes_core/sb1 [20]), .B(
        \U1/aes_core/sb0 [28]), .Y(\U1/aes_core/MC0/n33 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U93  ( .A(\U1/aes_core/MC0/n74 ), .B(
        \U1/aes_core/MC0/n33 ), .Y(\U1/aes_core/MC0/n20 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U92  ( .A(\U1/aes_core/MC0/n20 ), .B(
        \U1/aes_core/sb3 [4]), .Y(\U1/aes_core/MC0/n73 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U91  ( .A(\U1/aes_core/MC0/n54 ), .B(
        \U1/aes_core/MC0/n73 ), .Y(\U1/aes_core/sc0 [12]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U90  ( .A(\U1/aes_core/sb2 [12]), .B(
        \U1/aes_core/sb3 [4]), .Y(\U1/aes_core/MC0/n57 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U89  ( .A(\U1/aes_core/sb1 [21]), .B(
        \U1/aes_core/sb0 [29]), .Y(\U1/aes_core/MC0/n17 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U88  ( .A(\U1/aes_core/sb3 [5]), .B(
        \U1/aes_core/MC0/n17 ), .Y(\U1/aes_core/MC0/n72 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U87  ( .A(\U1/aes_core/MC0/n57 ), .B(
        \U1/aes_core/MC0/n72 ), .Y(\U1/aes_core/sc0 [13]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U86  ( .A(\U1/aes_core/sb2 [13]), .B(
        \U1/aes_core/sb3 [5]), .Y(\U1/aes_core/MC0/n31 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U85  ( .A(\U1/aes_core/sb1 [22]), .B(
        \U1/aes_core/sb0 [30]), .Y(\U1/aes_core/MC0/n14 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U84  ( .A(\U1/aes_core/sb3 [6]), .B(
        \U1/aes_core/MC0/n14 ), .Y(\U1/aes_core/MC0/n71 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U83  ( .A(\U1/aes_core/MC0/n31 ), .B(
        \U1/aes_core/MC0/n71 ), .Y(\U1/aes_core/sc0 [14]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U82  ( .A(\U1/aes_core/MC0/n11 ), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/MC0/n49 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U81  ( .A(\U1/aes_core/sb2 [14]), .B(
        \U1/aes_core/sb3 [6]), .Y(\U1/aes_core/MC0/n26 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U80  ( .A(\U1/aes_core/sb1 [23]), .B(
        \U1/aes_core/MC0/n26 ), .Y(\U1/aes_core/MC0/n70 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U79  ( .A(\U1/aes_core/MC0/n49 ), .B(
        \U1/aes_core/MC0/n70 ), .Y(\U1/aes_core/sc0 [15]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U78  ( .A(\U1/aes_core/sb0 [24]), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/MC0/n5 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U77  ( .A(\U1/aes_core/sb2 [8]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/MC0/n69 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U76  ( .A(\U1/aes_core/MC0/n69 ), .B(
        \U1/aes_core/sb3 [0]), .Y(\U1/aes_core/MC0/n45 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U75  ( .A(\U1/aes_core/MC0/n5 ), .B(
        \U1/aes_core/MC0/n45 ), .Y(\U1/aes_core/sc0 [16]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U74  ( .A(\U1/aes_core/sb1 [16]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/MC0/n67 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U73  ( .A(\U1/aes_core/MC0/n67 ), .B(
        \U1/aes_core/MC0/n68 ), .Y(\U1/aes_core/MC0/n44 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U72  ( .A(\U1/aes_core/MC0/n66 ), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/MC0/n3 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U71  ( .A(\U1/aes_core/sb0 [25]), .B(
        \U1/aes_core/MC0/n3 ), .Y(\U1/aes_core/MC0/n65 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U70  ( .A(\U1/aes_core/MC0/n44 ), .B(
        \U1/aes_core/MC0/n65 ), .Y(\U1/aes_core/sc0 [17]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U69  ( .A(\U1/aes_core/sb2 [9]), .B(
        \U1/aes_core/sb1 [17]), .Y(\U1/aes_core/MC0/n62 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U68  ( .A(\U1/aes_core/sb2 [10]), .B(
        \U1/aes_core/MC0/n64 ), .Y(\U1/aes_core/MC0/n63 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U67  ( .A(\U1/aes_core/MC0/n62 ), .B(
        \U1/aes_core/MC0/n63 ), .Y(\U1/aes_core/sc0 [18]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U66  ( .A(\U1/aes_core/sb2 [11]), .B(
        \U1/aes_core/sb1 [18]), .Y(\U1/aes_core/MC0/n60 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U65  ( .A(\U1/aes_core/sb3 [3]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/MC0/n61 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U64  ( .A(\U1/aes_core/MC0/n60 ), .B(
        \U1/aes_core/MC0/n61 ), .Y(\U1/aes_core/MC0/n38 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U63  ( .A(\U1/aes_core/MC0/n38 ), .B(
        \U1/aes_core/MC0/n59 ), .Y(\U1/aes_core/sc0 [19]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U62  ( .A(\U1/aes_core/sb0 [24]), .B(
        \U1/aes_core/sb0 [31]), .Y(\U1/aes_core/MC0/n42 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U61  ( .A(\U1/aes_core/sb1 [17]), .B(
        \U1/aes_core/sb0 [25]), .Y(\U1/aes_core/MC0/n41 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U60  ( .A(\U1/aes_core/sb3 [0]), .B(
        \U1/aes_core/sb3 [7]), .Y(\U1/aes_core/MC0/n7 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U59  ( .A(\U1/aes_core/MC0/n41 ), .B(
        \U1/aes_core/MC0/n7 ), .Y(\U1/aes_core/MC0/n4 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U58  ( .A(\U1/aes_core/MC0/n4 ), .B(
        \U1/aes_core/sb2 [9]), .Y(\U1/aes_core/MC0/n58 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U57  ( .A(\U1/aes_core/MC0/n42 ), .B(
        \U1/aes_core/MC0/n58 ), .Y(\U1/aes_core/sc0 [1]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U56  ( .A(\U1/aes_core/sb1 [19]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/MC0/n56 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U55  ( .A(\U1/aes_core/MC0/n56 ), .B(
        \U1/aes_core/MC0/n57 ), .Y(\U1/aes_core/MC0/n36 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U54  ( .A(\U1/aes_core/MC0/n36 ), .B(
        \U1/aes_core/sb0 [28]), .Y(\U1/aes_core/MC0/n55 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U53  ( .A(\U1/aes_core/MC0/n54 ), .B(
        \U1/aes_core/MC0/n55 ), .Y(\U1/aes_core/sc0 [20]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U52  ( .A(\U1/aes_core/sb0 [29]), .B(
        \U1/aes_core/sb1 [20]), .Y(\U1/aes_core/MC0/n52 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U51  ( .A(\U1/aes_core/sb2 [12]), .B(
        \U1/aes_core/MC0/n31 ), .Y(\U1/aes_core/MC0/n53 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U50  ( .A(\U1/aes_core/MC0/n52 ), .B(
        \U1/aes_core/MC0/n53 ), .Y(\U1/aes_core/sc0 [21]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U49  ( .A(\U1/aes_core/sb0 [30]), .B(
        \U1/aes_core/sb1 [21]), .Y(\U1/aes_core/MC0/n50 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U48  ( .A(\U1/aes_core/sb2 [13]), .B(
        \U1/aes_core/MC0/n26 ), .Y(\U1/aes_core/MC0/n51 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U47  ( .A(\U1/aes_core/MC0/n50 ), .B(
        \U1/aes_core/MC0/n51 ), .Y(\U1/aes_core/sc0 [22]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U46  ( .A(\U1/aes_core/sb1 [22]), .B(
        \U1/aes_core/sb2 [15]), .Y(\U1/aes_core/MC0/n47 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U45  ( .A(\U1/aes_core/sb2 [14]), .B(
        \U1/aes_core/MC0/n49 ), .Y(\U1/aes_core/MC0/n48 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U44  ( .A(\U1/aes_core/MC0/n47 ), .B(
        \U1/aes_core/MC0/n48 ), .Y(\U1/aes_core/sc0 [23]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U43  ( .A(\U1/aes_core/MC0/n45 ), .B(
        \U1/aes_core/MC0/n46 ), .Y(\U1/aes_core/sc0 [24]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U42  ( .A(\U1/aes_core/MC0/n44 ), .B(
        \U1/aes_core/sb1 [17]), .Y(\U1/aes_core/MC0/n43 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U41  ( .A(\U1/aes_core/MC0/n42 ), .B(
        \U1/aes_core/MC0/n43 ), .Y(\U1/aes_core/sc0 [25]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U40  ( .A(\U1/aes_core/sb2 [10]), .B(
        \U1/aes_core/sb1 [18]), .Y(\U1/aes_core/MC0/n30 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U39  ( .A(\U1/aes_core/sb3 [2]), .B(
        \U1/aes_core/MC0/n41 ), .Y(\U1/aes_core/MC0/n40 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U38  ( .A(\U1/aes_core/MC0/n30 ), .B(
        \U1/aes_core/MC0/n40 ), .Y(\U1/aes_core/sc0 [26]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U37  ( .A(\U1/aes_core/sb0 [26]), .B(
        \U1/aes_core/sb0 [31]), .Y(\U1/aes_core/MC0/n39 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U36  ( .A(\U1/aes_core/MC0/n39 ), .B(
        \U1/aes_core/sb1 [19]), .Y(\U1/aes_core/MC0/n23 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U32  ( .A(\U1/aes_core/sb0 [27]), .B(
        \U1/aes_core/MC0/n11 ), .Y(\U1/aes_core/MC0/n18 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U31  ( .A(\U1/aes_core/sb1 [20]), .B(
        \U1/aes_core/MC0/n18 ), .Y(\U1/aes_core/MC0/n35 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U29  ( .A(\U1/aes_core/sb1 [21]), .B(
        \U1/aes_core/MC0/n33 ), .Y(\U1/aes_core/MC0/n32 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U28  ( .A(\U1/aes_core/MC0/n31 ), .B(
        \U1/aes_core/MC0/n32 ), .Y(\U1/aes_core/sc0 [29]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U27  ( .A(\U1/aes_core/sb0 [26]), .B(
        \U1/aes_core/sb0 [25]), .Y(\U1/aes_core/MC0/n28 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U26  ( .A(\U1/aes_core/sb3 [1]), .B(
        \U1/aes_core/MC0/n30 ), .Y(\U1/aes_core/MC0/n29 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U25  ( .A(\U1/aes_core/MC0/n28 ), .B(
        \U1/aes_core/MC0/n29 ), .Y(\U1/aes_core/sc0 [2]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U24  ( .A(\U1/aes_core/sb1 [22]), .B(
        \U1/aes_core/MC0/n17 ), .Y(\U1/aes_core/MC0/n27 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U23  ( .A(\U1/aes_core/MC0/n26 ), .B(
        \U1/aes_core/MC0/n27 ), .Y(\U1/aes_core/sc0 [30]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U22  ( .A(\U1/aes_core/sb2 [15]), .B(
        \U1/aes_core/sb1 [23]), .Y(\U1/aes_core/MC0/n10 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U21  ( .A(\U1/aes_core/sb3 [7]), .B(
        \U1/aes_core/MC0/n10 ), .Y(\U1/aes_core/MC0/n25 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U20  ( .A(\U1/aes_core/MC0/n14 ), .B(
        \U1/aes_core/MC0/n25 ), .Y(\U1/aes_core/sc0 [31]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U19  ( .A(\U1/aes_core/sb2 [11]), .B(
        \U1/aes_core/sb0 [27]), .Y(\U1/aes_core/MC0/n21 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U18  ( .A(\U1/aes_core/MC0/n23 ), .B(
        \U1/aes_core/MC0/n24 ), .Y(\U1/aes_core/MC0/n22 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U17  ( .A(\U1/aes_core/MC0/n21 ), .B(
        \U1/aes_core/MC0/n22 ), .Y(\U1/aes_core/sc0 [3]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U16  ( .A(\U1/aes_core/MC0/n20 ), .B(
        \U1/aes_core/sb2 [12]), .Y(\U1/aes_core/MC0/n19 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U15  ( .A(\U1/aes_core/MC0/n18 ), .B(
        \U1/aes_core/MC0/n19 ), .Y(\U1/aes_core/sc0 [4]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U14  ( .A(\U1/aes_core/sb3 [4]), .B(
        \U1/aes_core/sb0 [28]), .Y(\U1/aes_core/MC0/n15 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U13  ( .A(\U1/aes_core/sb2 [13]), .B(
        \U1/aes_core/MC0/n17 ), .Y(\U1/aes_core/MC0/n16 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U12  ( .A(\U1/aes_core/MC0/n15 ), .B(
        \U1/aes_core/MC0/n16 ), .Y(\U1/aes_core/sc0 [5]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U11  ( .A(\U1/aes_core/sb3 [5]), .B(
        \U1/aes_core/sb0 [29]), .Y(\U1/aes_core/MC0/n12 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U10  ( .A(\U1/aes_core/sb2 [14]), .B(
        \U1/aes_core/MC0/n14 ), .Y(\U1/aes_core/MC0/n13 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U9  ( .A(\U1/aes_core/MC0/n12 ), .B(
        \U1/aes_core/MC0/n13 ), .Y(\U1/aes_core/sc0 [6]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC0/U8  ( .A(\U1/aes_core/sb3 [6]), .B(
        \U1/aes_core/MC0/n11 ), .Y(\U1/aes_core/MC0/n8 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U7  ( .A(\U1/aes_core/sb0 [30]), .B(
        \U1/aes_core/MC0/n10 ), .Y(\U1/aes_core/MC0/n9 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U6  ( .A(\U1/aes_core/MC0/n8 ), .B(
        \U1/aes_core/MC0/n9 ), .Y(\U1/aes_core/sc0 [7]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U5  ( .A(\U1/aes_core/sb1 [16]), .B(
        \U1/aes_core/MC0/n7 ), .Y(\U1/aes_core/MC0/n6 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U4  ( .A(\U1/aes_core/MC0/n5 ), .B(
        \U1/aes_core/MC0/n6 ), .Y(\U1/aes_core/sc0 [8]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC0/U2  ( .A(\U1/aes_core/sb3 [1]), .B(
        \U1/aes_core/MC0/n3 ), .Y(\U1/aes_core/MC0/n2 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U30  ( .A(\U1/aes_core/MC1/n118 ), .B(
        \U1/aes_core/MC1/n119 ), .Y(\U1/aes_core/sc1 [28]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U3  ( .A(\U1/aes_core/MC1/n130 ), .B(
        \U1/aes_core/MC1/n117 ), .Y(\U1/aes_core/sc1 [27]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U1  ( .A(\U1/aes_core/MC1/n149 ), .B(
        \U1/aes_core/MC1/n151 ), .Y(\U1/aes_core/sc1 [9]) );
  INV_X0P5B_A12TL \U1/aes_core/MC1/U112  ( .A(\U1/aes_core/sb3 [8]), .Y(
        \U1/aes_core/MC1/n89 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U111  ( .A(\U1/aes_core/MC1/n89 ), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/MC1/n34 ) );
  INV_X0P5B_A12TL \U1/aes_core/MC1/U110  ( .A(\U1/aes_core/sb1 [31]), .Y(
        \U1/aes_core/MC1/n142 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U109  ( .A(\U1/aes_core/sb2 [16]), .B(
        \U1/aes_core/MC1/n142 ), .Y(\U1/aes_core/MC1/n109 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U108  ( .A(\U1/aes_core/sb1 [24]), .B(
        \U1/aes_core/MC1/n109 ), .Y(\U1/aes_core/MC1/n1 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U107  ( .A(\U1/aes_core/MC1/n34 ), .B(
        \U1/aes_core/MC1/n1 ), .Y(\U1/aes_core/sc1 [0]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U106  ( .A(\U1/aes_core/sb1 [26]), .B(
        \U1/aes_core/sb0 [2]), .Y(\U1/aes_core/MC1/n91 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U105  ( .A(\U1/aes_core/sb0 [1]), .B(
        \U1/aes_core/sb3 [9]), .Y(\U1/aes_core/MC1/n87 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U104  ( .A(\U1/aes_core/sb2 [18]), .B(
        \U1/aes_core/MC1/n87 ), .Y(\U1/aes_core/MC1/n37 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U103  ( .A(\U1/aes_core/MC1/n91 ), .B(
        \U1/aes_core/MC1/n37 ), .Y(\U1/aes_core/sc1 [10]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U102  ( .A(\U1/aes_core/sb2 [19]), .B(
        \U1/aes_core/sb0 [3]), .Y(\U1/aes_core/MC1/n80 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U101  ( .A(\U1/aes_core/sb1 [27]), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/MC1/n78 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U100  ( .A(\U1/aes_core/MC1/n78 ), .B(
        \U1/aes_core/sb3 [10]), .Y(\U1/aes_core/MC1/n96 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U99  ( .A(\U1/aes_core/sb0 [2]), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/MC1/n129 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U98  ( .A(\U1/aes_core/MC1/n96 ), .B(
        \U1/aes_core/MC1/n129 ), .Y(\U1/aes_core/MC1/n79 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U97  ( .A(\U1/aes_core/MC1/n80 ), .B(
        \U1/aes_core/MC1/n79 ), .Y(\U1/aes_core/sc1 [11]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U96  ( .A(\U1/aes_core/sb3 [11]), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/MC1/n101 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U95  ( .A(\U1/aes_core/sb0 [3]), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/MC1/n81 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U94  ( .A(\U1/aes_core/sb2 [20]), .B(
        \U1/aes_core/sb1 [28]), .Y(\U1/aes_core/MC1/n120 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U93  ( .A(\U1/aes_core/MC1/n81 ), .B(
        \U1/aes_core/MC1/n120 ), .Y(\U1/aes_core/MC1/n133 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U92  ( .A(\U1/aes_core/MC1/n133 ), .B(
        \U1/aes_core/sb0 [4]), .Y(\U1/aes_core/MC1/n82 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U91  ( .A(\U1/aes_core/MC1/n101 ), .B(
        \U1/aes_core/MC1/n82 ), .Y(\U1/aes_core/sc1 [12]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U90  ( .A(\U1/aes_core/sb3 [12]), .B(
        \U1/aes_core/sb0 [4]), .Y(\U1/aes_core/MC1/n98 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U89  ( .A(\U1/aes_core/sb2 [21]), .B(
        \U1/aes_core/sb1 [29]), .Y(\U1/aes_core/MC1/n136 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U88  ( .A(\U1/aes_core/sb0 [5]), .B(
        \U1/aes_core/MC1/n136 ), .Y(\U1/aes_core/MC1/n83 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U87  ( .A(\U1/aes_core/MC1/n98 ), .B(
        \U1/aes_core/MC1/n83 ), .Y(\U1/aes_core/sc1 [13]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U86  ( .A(\U1/aes_core/sb3 [13]), .B(
        \U1/aes_core/sb0 [5]), .Y(\U1/aes_core/MC1/n122 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U85  ( .A(\U1/aes_core/sb2 [22]), .B(
        \U1/aes_core/sb1 [30]), .Y(\U1/aes_core/MC1/n139 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U84  ( .A(\U1/aes_core/sb0 [6]), .B(
        \U1/aes_core/MC1/n139 ), .Y(\U1/aes_core/MC1/n84 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U83  ( .A(\U1/aes_core/MC1/n122 ), .B(
        \U1/aes_core/MC1/n84 ), .Y(\U1/aes_core/sc1 [14]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U82  ( .A(\U1/aes_core/MC1/n142 ), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/MC1/n106 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U81  ( .A(\U1/aes_core/sb3 [14]), .B(
        \U1/aes_core/sb0 [6]), .Y(\U1/aes_core/MC1/n127 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U80  ( .A(\U1/aes_core/sb2 [23]), .B(
        \U1/aes_core/MC1/n127 ), .Y(\U1/aes_core/MC1/n85 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U79  ( .A(\U1/aes_core/MC1/n106 ), .B(
        \U1/aes_core/MC1/n85 ), .Y(\U1/aes_core/sc1 [15]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U78  ( .A(\U1/aes_core/sb1 [24]), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/MC1/n148 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U77  ( .A(\U1/aes_core/sb3 [8]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/MC1/n86 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U76  ( .A(\U1/aes_core/MC1/n86 ), .B(
        \U1/aes_core/sb0 [0]), .Y(\U1/aes_core/MC1/n110 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U75  ( .A(\U1/aes_core/MC1/n148 ), .B(
        \U1/aes_core/MC1/n110 ), .Y(\U1/aes_core/sc1 [16]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U74  ( .A(\U1/aes_core/sb2 [16]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/MC1/n88 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U73  ( .A(\U1/aes_core/MC1/n88 ), .B(
        \U1/aes_core/MC1/n87 ), .Y(\U1/aes_core/MC1/n111 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U72  ( .A(\U1/aes_core/MC1/n89 ), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/MC1/n150 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U71  ( .A(\U1/aes_core/sb1 [25]), .B(
        \U1/aes_core/MC1/n150 ), .Y(\U1/aes_core/MC1/n90 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U70  ( .A(\U1/aes_core/MC1/n111 ), .B(
        \U1/aes_core/MC1/n90 ), .Y(\U1/aes_core/sc1 [17]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U69  ( .A(\U1/aes_core/sb3 [9]), .B(
        \U1/aes_core/sb2 [17]), .Y(\U1/aes_core/MC1/n93 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U68  ( .A(\U1/aes_core/sb3 [10]), .B(
        \U1/aes_core/MC1/n91 ), .Y(\U1/aes_core/MC1/n92 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U67  ( .A(\U1/aes_core/MC1/n93 ), .B(
        \U1/aes_core/MC1/n92 ), .Y(\U1/aes_core/sc1 [18]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U66  ( .A(\U1/aes_core/sb3 [11]), .B(
        \U1/aes_core/sb2 [18]), .Y(\U1/aes_core/MC1/n95 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U65  ( .A(\U1/aes_core/sb0 [3]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/MC1/n94 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U64  ( .A(\U1/aes_core/MC1/n95 ), .B(
        \U1/aes_core/MC1/n94 ), .Y(\U1/aes_core/MC1/n117 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U63  ( .A(\U1/aes_core/MC1/n117 ), .B(
        \U1/aes_core/MC1/n96 ), .Y(\U1/aes_core/sc1 [19]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U62  ( .A(\U1/aes_core/sb1 [24]), .B(
        \U1/aes_core/sb1 [31]), .Y(\U1/aes_core/MC1/n113 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U61  ( .A(\U1/aes_core/sb2 [17]), .B(
        \U1/aes_core/sb1 [25]), .Y(\U1/aes_core/MC1/n114 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U60  ( .A(\U1/aes_core/sb0 [0]), .B(
        \U1/aes_core/sb0 [7]), .Y(\U1/aes_core/MC1/n146 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U59  ( .A(\U1/aes_core/MC1/n114 ), .B(
        \U1/aes_core/MC1/n146 ), .Y(\U1/aes_core/MC1/n149 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U58  ( .A(\U1/aes_core/MC1/n149 ), .B(
        \U1/aes_core/sb3 [9]), .Y(\U1/aes_core/MC1/n97 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U57  ( .A(\U1/aes_core/MC1/n113 ), .B(
        \U1/aes_core/MC1/n97 ), .Y(\U1/aes_core/sc1 [1]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U56  ( .A(\U1/aes_core/sb2 [19]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/MC1/n99 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U55  ( .A(\U1/aes_core/MC1/n99 ), .B(
        \U1/aes_core/MC1/n98 ), .Y(\U1/aes_core/MC1/n118 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U54  ( .A(\U1/aes_core/MC1/n118 ), .B(
        \U1/aes_core/sb1 [28]), .Y(\U1/aes_core/MC1/n100 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U53  ( .A(\U1/aes_core/MC1/n101 ), .B(
        \U1/aes_core/MC1/n100 ), .Y(\U1/aes_core/sc1 [20]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U52  ( .A(\U1/aes_core/sb1 [29]), .B(
        \U1/aes_core/sb2 [20]), .Y(\U1/aes_core/MC1/n103 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U51  ( .A(\U1/aes_core/sb3 [12]), .B(
        \U1/aes_core/MC1/n122 ), .Y(\U1/aes_core/MC1/n102 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U50  ( .A(\U1/aes_core/MC1/n103 ), .B(
        \U1/aes_core/MC1/n102 ), .Y(\U1/aes_core/sc1 [21]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U49  ( .A(\U1/aes_core/sb1 [30]), .B(
        \U1/aes_core/sb2 [21]), .Y(\U1/aes_core/MC1/n105 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U48  ( .A(\U1/aes_core/sb3 [13]), .B(
        \U1/aes_core/MC1/n127 ), .Y(\U1/aes_core/MC1/n104 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U47  ( .A(\U1/aes_core/MC1/n105 ), .B(
        \U1/aes_core/MC1/n104 ), .Y(\U1/aes_core/sc1 [22]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U46  ( .A(\U1/aes_core/sb2 [22]), .B(
        \U1/aes_core/sb3 [15]), .Y(\U1/aes_core/MC1/n108 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U45  ( .A(\U1/aes_core/sb3 [14]), .B(
        \U1/aes_core/MC1/n106 ), .Y(\U1/aes_core/MC1/n107 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U44  ( .A(\U1/aes_core/MC1/n108 ), .B(
        \U1/aes_core/MC1/n107 ), .Y(\U1/aes_core/sc1 [23]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U43  ( .A(\U1/aes_core/MC1/n110 ), .B(
        \U1/aes_core/MC1/n109 ), .Y(\U1/aes_core/sc1 [24]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U42  ( .A(\U1/aes_core/MC1/n111 ), .B(
        \U1/aes_core/sb2 [17]), .Y(\U1/aes_core/MC1/n112 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U41  ( .A(\U1/aes_core/MC1/n113 ), .B(
        \U1/aes_core/MC1/n112 ), .Y(\U1/aes_core/sc1 [25]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U40  ( .A(\U1/aes_core/sb3 [10]), .B(
        \U1/aes_core/sb2 [18]), .Y(\U1/aes_core/MC1/n123 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U39  ( .A(\U1/aes_core/sb0 [2]), .B(
        \U1/aes_core/MC1/n114 ), .Y(\U1/aes_core/MC1/n115 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U38  ( .A(\U1/aes_core/MC1/n123 ), .B(
        \U1/aes_core/MC1/n115 ), .Y(\U1/aes_core/sc1 [26]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U37  ( .A(\U1/aes_core/sb1 [26]), .B(
        \U1/aes_core/sb1 [31]), .Y(\U1/aes_core/MC1/n116 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U36  ( .A(\U1/aes_core/MC1/n116 ), .B(
        \U1/aes_core/sb2 [19]), .Y(\U1/aes_core/MC1/n130 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U32  ( .A(\U1/aes_core/sb1 [27]), .B(
        \U1/aes_core/MC1/n142 ), .Y(\U1/aes_core/MC1/n135 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U31  ( .A(\U1/aes_core/sb2 [20]), .B(
        \U1/aes_core/MC1/n135 ), .Y(\U1/aes_core/MC1/n119 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U29  ( .A(\U1/aes_core/sb2 [21]), .B(
        \U1/aes_core/MC1/n120 ), .Y(\U1/aes_core/MC1/n121 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U28  ( .A(\U1/aes_core/MC1/n122 ), .B(
        \U1/aes_core/MC1/n121 ), .Y(\U1/aes_core/sc1 [29]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U27  ( .A(\U1/aes_core/sb1 [26]), .B(
        \U1/aes_core/sb1 [25]), .Y(\U1/aes_core/MC1/n125 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U26  ( .A(\U1/aes_core/sb0 [1]), .B(
        \U1/aes_core/MC1/n123 ), .Y(\U1/aes_core/MC1/n124 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U25  ( .A(\U1/aes_core/MC1/n125 ), .B(
        \U1/aes_core/MC1/n124 ), .Y(\U1/aes_core/sc1 [2]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U24  ( .A(\U1/aes_core/sb2 [22]), .B(
        \U1/aes_core/MC1/n136 ), .Y(\U1/aes_core/MC1/n126 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U23  ( .A(\U1/aes_core/MC1/n127 ), .B(
        \U1/aes_core/MC1/n126 ), .Y(\U1/aes_core/sc1 [30]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U22  ( .A(\U1/aes_core/sb3 [15]), .B(
        \U1/aes_core/sb2 [23]), .Y(\U1/aes_core/MC1/n143 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U21  ( .A(\U1/aes_core/sb0 [7]), .B(
        \U1/aes_core/MC1/n143 ), .Y(\U1/aes_core/MC1/n128 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U20  ( .A(\U1/aes_core/MC1/n139 ), .B(
        \U1/aes_core/MC1/n128 ), .Y(\U1/aes_core/sc1 [31]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U19  ( .A(\U1/aes_core/sb3 [11]), .B(
        \U1/aes_core/sb1 [27]), .Y(\U1/aes_core/MC1/n132 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U18  ( .A(\U1/aes_core/MC1/n130 ), .B(
        \U1/aes_core/MC1/n129 ), .Y(\U1/aes_core/MC1/n131 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U17  ( .A(\U1/aes_core/MC1/n132 ), .B(
        \U1/aes_core/MC1/n131 ), .Y(\U1/aes_core/sc1 [3]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U16  ( .A(\U1/aes_core/MC1/n133 ), .B(
        \U1/aes_core/sb3 [12]), .Y(\U1/aes_core/MC1/n134 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U15  ( .A(\U1/aes_core/MC1/n135 ), .B(
        \U1/aes_core/MC1/n134 ), .Y(\U1/aes_core/sc1 [4]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U14  ( .A(\U1/aes_core/sb0 [4]), .B(
        \U1/aes_core/sb1 [28]), .Y(\U1/aes_core/MC1/n138 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U13  ( .A(\U1/aes_core/sb3 [13]), .B(
        \U1/aes_core/MC1/n136 ), .Y(\U1/aes_core/MC1/n137 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U12  ( .A(\U1/aes_core/MC1/n138 ), .B(
        \U1/aes_core/MC1/n137 ), .Y(\U1/aes_core/sc1 [5]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U11  ( .A(\U1/aes_core/sb0 [5]), .B(
        \U1/aes_core/sb1 [29]), .Y(\U1/aes_core/MC1/n141 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U10  ( .A(\U1/aes_core/sb3 [14]), .B(
        \U1/aes_core/MC1/n139 ), .Y(\U1/aes_core/MC1/n140 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U9  ( .A(\U1/aes_core/MC1/n141 ), .B(
        \U1/aes_core/MC1/n140 ), .Y(\U1/aes_core/sc1 [6]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC1/U8  ( .A(\U1/aes_core/sb0 [6]), .B(
        \U1/aes_core/MC1/n142 ), .Y(\U1/aes_core/MC1/n145 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U7  ( .A(\U1/aes_core/sb1 [30]), .B(
        \U1/aes_core/MC1/n143 ), .Y(\U1/aes_core/MC1/n144 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U6  ( .A(\U1/aes_core/MC1/n145 ), .B(
        \U1/aes_core/MC1/n144 ), .Y(\U1/aes_core/sc1 [7]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U5  ( .A(\U1/aes_core/sb2 [16]), .B(
        \U1/aes_core/MC1/n146 ), .Y(\U1/aes_core/MC1/n147 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U4  ( .A(\U1/aes_core/MC1/n148 ), .B(
        \U1/aes_core/MC1/n147 ), .Y(\U1/aes_core/sc1 [8]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC1/U2  ( .A(\U1/aes_core/sb0 [1]), .B(
        \U1/aes_core/MC1/n150 ), .Y(\U1/aes_core/MC1/n151 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U30  ( .A(\U1/aes_core/MC2/n118 ), .B(
        \U1/aes_core/MC2/n119 ), .Y(\U1/aes_core/sc2 [28]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U3  ( .A(\U1/aes_core/MC2/n130 ), .B(
        \U1/aes_core/MC2/n117 ), .Y(\U1/aes_core/sc2 [27]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U1  ( .A(\U1/aes_core/MC2/n149 ), .B(
        \U1/aes_core/MC2/n151 ), .Y(\U1/aes_core/sc2 [9]) );
  INV_X0P5B_A12TL \U1/aes_core/MC2/U112  ( .A(\U1/aes_core/sb0 [8]), .Y(
        \U1/aes_core/MC2/n89 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U111  ( .A(\U1/aes_core/MC2/n89 ), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/MC2/n34 ) );
  INV_X0P5B_A12TL \U1/aes_core/MC2/U110  ( .A(\U1/aes_core/sb2 [31]), .Y(
        \U1/aes_core/MC2/n142 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U109  ( .A(\U1/aes_core/sb3 [16]), .B(
        \U1/aes_core/MC2/n142 ), .Y(\U1/aes_core/MC2/n109 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U108  ( .A(\U1/aes_core/sb2 [24]), .B(
        \U1/aes_core/MC2/n109 ), .Y(\U1/aes_core/MC2/n1 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U107  ( .A(\U1/aes_core/MC2/n34 ), .B(
        \U1/aes_core/MC2/n1 ), .Y(\U1/aes_core/sc2 [0]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U106  ( .A(\U1/aes_core/sb2 [26]), .B(
        \U1/aes_core/sb1 [2]), .Y(\U1/aes_core/MC2/n91 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U105  ( .A(\U1/aes_core/sb1 [1]), .B(
        \U1/aes_core/sb0 [9]), .Y(\U1/aes_core/MC2/n87 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U104  ( .A(\U1/aes_core/sb3 [18]), .B(
        \U1/aes_core/MC2/n87 ), .Y(\U1/aes_core/MC2/n37 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U103  ( .A(\U1/aes_core/MC2/n91 ), .B(
        \U1/aes_core/MC2/n37 ), .Y(\U1/aes_core/sc2 [10]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U102  ( .A(\U1/aes_core/sb3 [19]), .B(
        \U1/aes_core/sb1 [3]), .Y(\U1/aes_core/MC2/n80 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U101  ( .A(\U1/aes_core/sb2 [27]), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/MC2/n78 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U100  ( .A(\U1/aes_core/MC2/n78 ), .B(
        \U1/aes_core/sb0 [10]), .Y(\U1/aes_core/MC2/n96 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U99  ( .A(\U1/aes_core/sb1 [2]), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/MC2/n129 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U98  ( .A(\U1/aes_core/MC2/n96 ), .B(
        \U1/aes_core/MC2/n129 ), .Y(\U1/aes_core/MC2/n79 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U97  ( .A(\U1/aes_core/MC2/n80 ), .B(
        \U1/aes_core/MC2/n79 ), .Y(\U1/aes_core/sc2 [11]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U96  ( .A(\U1/aes_core/sb0 [11]), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/MC2/n101 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U95  ( .A(\U1/aes_core/sb1 [3]), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/MC2/n81 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U94  ( .A(\U1/aes_core/sb3 [20]), .B(
        \U1/aes_core/sb2 [28]), .Y(\U1/aes_core/MC2/n120 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U93  ( .A(\U1/aes_core/MC2/n81 ), .B(
        \U1/aes_core/MC2/n120 ), .Y(\U1/aes_core/MC2/n133 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U92  ( .A(\U1/aes_core/MC2/n133 ), .B(
        \U1/aes_core/sb1 [4]), .Y(\U1/aes_core/MC2/n82 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U91  ( .A(\U1/aes_core/MC2/n101 ), .B(
        \U1/aes_core/MC2/n82 ), .Y(\U1/aes_core/sc2 [12]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U90  ( .A(\U1/aes_core/sb0 [12]), .B(
        \U1/aes_core/sb1 [4]), .Y(\U1/aes_core/MC2/n98 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U89  ( .A(\U1/aes_core/sb3 [21]), .B(
        \U1/aes_core/sb2 [29]), .Y(\U1/aes_core/MC2/n136 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U88  ( .A(\U1/aes_core/sb1 [5]), .B(
        \U1/aes_core/MC2/n136 ), .Y(\U1/aes_core/MC2/n83 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U87  ( .A(\U1/aes_core/MC2/n98 ), .B(
        \U1/aes_core/MC2/n83 ), .Y(\U1/aes_core/sc2 [13]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U86  ( .A(\U1/aes_core/sb0 [13]), .B(
        \U1/aes_core/sb1 [5]), .Y(\U1/aes_core/MC2/n122 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U85  ( .A(\U1/aes_core/sb3 [22]), .B(
        \U1/aes_core/sb2 [30]), .Y(\U1/aes_core/MC2/n139 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U84  ( .A(\U1/aes_core/sb1 [6]), .B(
        \U1/aes_core/MC2/n139 ), .Y(\U1/aes_core/MC2/n84 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U83  ( .A(\U1/aes_core/MC2/n122 ), .B(
        \U1/aes_core/MC2/n84 ), .Y(\U1/aes_core/sc2 [14]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U82  ( .A(\U1/aes_core/MC2/n142 ), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/MC2/n106 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U81  ( .A(\U1/aes_core/sb0 [14]), .B(
        \U1/aes_core/sb1 [6]), .Y(\U1/aes_core/MC2/n127 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U80  ( .A(\U1/aes_core/sb3 [23]), .B(
        \U1/aes_core/MC2/n127 ), .Y(\U1/aes_core/MC2/n85 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U79  ( .A(\U1/aes_core/MC2/n106 ), .B(
        \U1/aes_core/MC2/n85 ), .Y(\U1/aes_core/sc2 [15]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U78  ( .A(\U1/aes_core/sb2 [24]), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/MC2/n148 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U77  ( .A(\U1/aes_core/sb0 [8]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/MC2/n86 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U76  ( .A(\U1/aes_core/MC2/n86 ), .B(
        \U1/aes_core/sb1 [0]), .Y(\U1/aes_core/MC2/n110 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U75  ( .A(\U1/aes_core/MC2/n148 ), .B(
        \U1/aes_core/MC2/n110 ), .Y(\U1/aes_core/sc2 [16]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U74  ( .A(\U1/aes_core/sb3 [16]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/MC2/n88 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U73  ( .A(\U1/aes_core/MC2/n88 ), .B(
        \U1/aes_core/MC2/n87 ), .Y(\U1/aes_core/MC2/n111 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U72  ( .A(\U1/aes_core/MC2/n89 ), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/MC2/n150 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U71  ( .A(\U1/aes_core/sb2 [25]), .B(
        \U1/aes_core/MC2/n150 ), .Y(\U1/aes_core/MC2/n90 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U70  ( .A(\U1/aes_core/MC2/n111 ), .B(
        \U1/aes_core/MC2/n90 ), .Y(\U1/aes_core/sc2 [17]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U69  ( .A(\U1/aes_core/sb0 [9]), .B(
        \U1/aes_core/sb3 [17]), .Y(\U1/aes_core/MC2/n93 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U68  ( .A(\U1/aes_core/sb0 [10]), .B(
        \U1/aes_core/MC2/n91 ), .Y(\U1/aes_core/MC2/n92 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U67  ( .A(\U1/aes_core/MC2/n93 ), .B(
        \U1/aes_core/MC2/n92 ), .Y(\U1/aes_core/sc2 [18]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U66  ( .A(\U1/aes_core/sb0 [11]), .B(
        \U1/aes_core/sb3 [18]), .Y(\U1/aes_core/MC2/n95 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U65  ( .A(\U1/aes_core/sb1 [3]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/MC2/n94 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U64  ( .A(\U1/aes_core/MC2/n95 ), .B(
        \U1/aes_core/MC2/n94 ), .Y(\U1/aes_core/MC2/n117 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U63  ( .A(\U1/aes_core/MC2/n117 ), .B(
        \U1/aes_core/MC2/n96 ), .Y(\U1/aes_core/sc2 [19]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U62  ( .A(\U1/aes_core/sb2 [24]), .B(
        \U1/aes_core/sb2 [31]), .Y(\U1/aes_core/MC2/n113 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U61  ( .A(\U1/aes_core/sb3 [17]), .B(
        \U1/aes_core/sb2 [25]), .Y(\U1/aes_core/MC2/n114 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U60  ( .A(\U1/aes_core/sb1 [0]), .B(
        \U1/aes_core/sb1 [7]), .Y(\U1/aes_core/MC2/n146 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U59  ( .A(\U1/aes_core/MC2/n114 ), .B(
        \U1/aes_core/MC2/n146 ), .Y(\U1/aes_core/MC2/n149 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U58  ( .A(\U1/aes_core/MC2/n149 ), .B(
        \U1/aes_core/sb0 [9]), .Y(\U1/aes_core/MC2/n97 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U57  ( .A(\U1/aes_core/MC2/n113 ), .B(
        \U1/aes_core/MC2/n97 ), .Y(\U1/aes_core/sc2 [1]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U56  ( .A(\U1/aes_core/sb3 [19]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/MC2/n99 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U55  ( .A(\U1/aes_core/MC2/n99 ), .B(
        \U1/aes_core/MC2/n98 ), .Y(\U1/aes_core/MC2/n118 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U54  ( .A(\U1/aes_core/MC2/n118 ), .B(
        \U1/aes_core/sb2 [28]), .Y(\U1/aes_core/MC2/n100 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U53  ( .A(\U1/aes_core/MC2/n101 ), .B(
        \U1/aes_core/MC2/n100 ), .Y(\U1/aes_core/sc2 [20]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U52  ( .A(\U1/aes_core/sb2 [29]), .B(
        \U1/aes_core/sb3 [20]), .Y(\U1/aes_core/MC2/n103 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U51  ( .A(\U1/aes_core/sb0 [12]), .B(
        \U1/aes_core/MC2/n122 ), .Y(\U1/aes_core/MC2/n102 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U50  ( .A(\U1/aes_core/MC2/n103 ), .B(
        \U1/aes_core/MC2/n102 ), .Y(\U1/aes_core/sc2 [21]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U49  ( .A(\U1/aes_core/sb2 [30]), .B(
        \U1/aes_core/sb3 [21]), .Y(\U1/aes_core/MC2/n105 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U48  ( .A(\U1/aes_core/sb0 [13]), .B(
        \U1/aes_core/MC2/n127 ), .Y(\U1/aes_core/MC2/n104 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U47  ( .A(\U1/aes_core/MC2/n105 ), .B(
        \U1/aes_core/MC2/n104 ), .Y(\U1/aes_core/sc2 [22]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U46  ( .A(\U1/aes_core/sb3 [22]), .B(
        \U1/aes_core/sb0 [15]), .Y(\U1/aes_core/MC2/n108 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U45  ( .A(\U1/aes_core/sb0 [14]), .B(
        \U1/aes_core/MC2/n106 ), .Y(\U1/aes_core/MC2/n107 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U44  ( .A(\U1/aes_core/MC2/n108 ), .B(
        \U1/aes_core/MC2/n107 ), .Y(\U1/aes_core/sc2 [23]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U43  ( .A(\U1/aes_core/MC2/n110 ), .B(
        \U1/aes_core/MC2/n109 ), .Y(\U1/aes_core/sc2 [24]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U42  ( .A(\U1/aes_core/MC2/n111 ), .B(
        \U1/aes_core/sb3 [17]), .Y(\U1/aes_core/MC2/n112 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U41  ( .A(\U1/aes_core/MC2/n113 ), .B(
        \U1/aes_core/MC2/n112 ), .Y(\U1/aes_core/sc2 [25]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U40  ( .A(\U1/aes_core/sb0 [10]), .B(
        \U1/aes_core/sb3 [18]), .Y(\U1/aes_core/MC2/n123 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U39  ( .A(\U1/aes_core/sb1 [2]), .B(
        \U1/aes_core/MC2/n114 ), .Y(\U1/aes_core/MC2/n115 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U38  ( .A(\U1/aes_core/MC2/n123 ), .B(
        \U1/aes_core/MC2/n115 ), .Y(\U1/aes_core/sc2 [26]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U37  ( .A(\U1/aes_core/sb2 [26]), .B(
        \U1/aes_core/sb2 [31]), .Y(\U1/aes_core/MC2/n116 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U36  ( .A(\U1/aes_core/MC2/n116 ), .B(
        \U1/aes_core/sb3 [19]), .Y(\U1/aes_core/MC2/n130 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U32  ( .A(\U1/aes_core/sb2 [27]), .B(
        \U1/aes_core/MC2/n142 ), .Y(\U1/aes_core/MC2/n135 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U31  ( .A(\U1/aes_core/sb3 [20]), .B(
        \U1/aes_core/MC2/n135 ), .Y(\U1/aes_core/MC2/n119 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U29  ( .A(\U1/aes_core/sb3 [21]), .B(
        \U1/aes_core/MC2/n120 ), .Y(\U1/aes_core/MC2/n121 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U28  ( .A(\U1/aes_core/MC2/n122 ), .B(
        \U1/aes_core/MC2/n121 ), .Y(\U1/aes_core/sc2 [29]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U27  ( .A(\U1/aes_core/sb2 [26]), .B(
        \U1/aes_core/sb2 [25]), .Y(\U1/aes_core/MC2/n125 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U26  ( .A(\U1/aes_core/sb1 [1]), .B(
        \U1/aes_core/MC2/n123 ), .Y(\U1/aes_core/MC2/n124 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U25  ( .A(\U1/aes_core/MC2/n125 ), .B(
        \U1/aes_core/MC2/n124 ), .Y(\U1/aes_core/sc2 [2]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U24  ( .A(\U1/aes_core/sb3 [22]), .B(
        \U1/aes_core/MC2/n136 ), .Y(\U1/aes_core/MC2/n126 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U23  ( .A(\U1/aes_core/MC2/n127 ), .B(
        \U1/aes_core/MC2/n126 ), .Y(\U1/aes_core/sc2 [30]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U22  ( .A(\U1/aes_core/sb0 [15]), .B(
        \U1/aes_core/sb3 [23]), .Y(\U1/aes_core/MC2/n143 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U21  ( .A(\U1/aes_core/sb1 [7]), .B(
        \U1/aes_core/MC2/n143 ), .Y(\U1/aes_core/MC2/n128 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U20  ( .A(\U1/aes_core/MC2/n139 ), .B(
        \U1/aes_core/MC2/n128 ), .Y(\U1/aes_core/sc2 [31]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U19  ( .A(\U1/aes_core/sb0 [11]), .B(
        \U1/aes_core/sb2 [27]), .Y(\U1/aes_core/MC2/n132 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U18  ( .A(\U1/aes_core/MC2/n130 ), .B(
        \U1/aes_core/MC2/n129 ), .Y(\U1/aes_core/MC2/n131 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U17  ( .A(\U1/aes_core/MC2/n132 ), .B(
        \U1/aes_core/MC2/n131 ), .Y(\U1/aes_core/sc2 [3]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U16  ( .A(\U1/aes_core/MC2/n133 ), .B(
        \U1/aes_core/sb0 [12]), .Y(\U1/aes_core/MC2/n134 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U15  ( .A(\U1/aes_core/MC2/n135 ), .B(
        \U1/aes_core/MC2/n134 ), .Y(\U1/aes_core/sc2 [4]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U14  ( .A(\U1/aes_core/sb1 [4]), .B(
        \U1/aes_core/sb2 [28]), .Y(\U1/aes_core/MC2/n138 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U13  ( .A(\U1/aes_core/sb0 [13]), .B(
        \U1/aes_core/MC2/n136 ), .Y(\U1/aes_core/MC2/n137 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U12  ( .A(\U1/aes_core/MC2/n138 ), .B(
        \U1/aes_core/MC2/n137 ), .Y(\U1/aes_core/sc2 [5]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U11  ( .A(\U1/aes_core/sb1 [5]), .B(
        \U1/aes_core/sb2 [29]), .Y(\U1/aes_core/MC2/n141 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U10  ( .A(\U1/aes_core/sb0 [14]), .B(
        \U1/aes_core/MC2/n139 ), .Y(\U1/aes_core/MC2/n140 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U9  ( .A(\U1/aes_core/MC2/n141 ), .B(
        \U1/aes_core/MC2/n140 ), .Y(\U1/aes_core/sc2 [6]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC2/U8  ( .A(\U1/aes_core/sb1 [6]), .B(
        \U1/aes_core/MC2/n142 ), .Y(\U1/aes_core/MC2/n145 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U7  ( .A(\U1/aes_core/sb2 [30]), .B(
        \U1/aes_core/MC2/n143 ), .Y(\U1/aes_core/MC2/n144 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U6  ( .A(\U1/aes_core/MC2/n145 ), .B(
        \U1/aes_core/MC2/n144 ), .Y(\U1/aes_core/sc2 [7]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U5  ( .A(\U1/aes_core/sb3 [16]), .B(
        \U1/aes_core/MC2/n146 ), .Y(\U1/aes_core/MC2/n147 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U4  ( .A(\U1/aes_core/MC2/n148 ), .B(
        \U1/aes_core/MC2/n147 ), .Y(\U1/aes_core/sc2 [8]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC2/U2  ( .A(\U1/aes_core/sb1 [1]), .B(
        \U1/aes_core/MC2/n150 ), .Y(\U1/aes_core/MC2/n151 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U30  ( .A(\U1/aes_core/MC3/n118 ), .B(
        \U1/aes_core/MC3/n119 ), .Y(\U1/aes_core/sc3 [28]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U3  ( .A(\U1/aes_core/MC3/n130 ), .B(
        \U1/aes_core/MC3/n117 ), .Y(\U1/aes_core/sc3 [27]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U1  ( .A(\U1/aes_core/MC3/n149 ), .B(
        \U1/aes_core/MC3/n151 ), .Y(\U1/aes_core/sc3 [9]) );
  INV_X0P5B_A12TL \U1/aes_core/MC3/U112  ( .A(\U1/aes_core/sb1 [8]), .Y(
        \U1/aes_core/MC3/n89 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U111  ( .A(\U1/aes_core/MC3/n89 ), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/MC3/n34 ) );
  INV_X0P5B_A12TL \U1/aes_core/MC3/U110  ( .A(\U1/aes_core/sb3 [31]), .Y(
        \U1/aes_core/MC3/n142 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U109  ( .A(\U1/aes_core/sb0 [16]), .B(
        \U1/aes_core/MC3/n142 ), .Y(\U1/aes_core/MC3/n109 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U108  ( .A(\U1/aes_core/sb3 [24]), .B(
        \U1/aes_core/MC3/n109 ), .Y(\U1/aes_core/MC3/n1 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U107  ( .A(\U1/aes_core/MC3/n34 ), .B(
        \U1/aes_core/MC3/n1 ), .Y(\U1/aes_core/sc3 [0]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U106  ( .A(\U1/aes_core/sb3 [26]), .B(
        \U1/aes_core/sb2 [2]), .Y(\U1/aes_core/MC3/n91 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U105  ( .A(\U1/aes_core/sb2 [1]), .B(
        \U1/aes_core/sb1 [9]), .Y(\U1/aes_core/MC3/n87 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U104  ( .A(\U1/aes_core/sb0 [18]), .B(
        \U1/aes_core/MC3/n87 ), .Y(\U1/aes_core/MC3/n37 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U103  ( .A(\U1/aes_core/MC3/n91 ), .B(
        \U1/aes_core/MC3/n37 ), .Y(\U1/aes_core/sc3 [10]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U102  ( .A(\U1/aes_core/sb0 [19]), .B(
        \U1/aes_core/sb2 [3]), .Y(\U1/aes_core/MC3/n80 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U101  ( .A(\U1/aes_core/sb3 [27]), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/MC3/n78 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U100  ( .A(\U1/aes_core/MC3/n78 ), .B(
        \U1/aes_core/sb1 [10]), .Y(\U1/aes_core/MC3/n96 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U99  ( .A(\U1/aes_core/sb2 [2]), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/MC3/n129 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U98  ( .A(\U1/aes_core/MC3/n96 ), .B(
        \U1/aes_core/MC3/n129 ), .Y(\U1/aes_core/MC3/n79 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U97  ( .A(\U1/aes_core/MC3/n80 ), .B(
        \U1/aes_core/MC3/n79 ), .Y(\U1/aes_core/sc3 [11]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U96  ( .A(\U1/aes_core/sb1 [11]), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/MC3/n101 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U95  ( .A(\U1/aes_core/sb2 [3]), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/MC3/n81 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U94  ( .A(\U1/aes_core/sb0 [20]), .B(
        \U1/aes_core/sb3 [28]), .Y(\U1/aes_core/MC3/n120 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U93  ( .A(\U1/aes_core/MC3/n81 ), .B(
        \U1/aes_core/MC3/n120 ), .Y(\U1/aes_core/MC3/n133 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U92  ( .A(\U1/aes_core/MC3/n133 ), .B(
        \U1/aes_core/sb2 [4]), .Y(\U1/aes_core/MC3/n82 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U91  ( .A(\U1/aes_core/MC3/n101 ), .B(
        \U1/aes_core/MC3/n82 ), .Y(\U1/aes_core/sc3 [12]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U90  ( .A(\U1/aes_core/sb1 [12]), .B(
        \U1/aes_core/sb2 [4]), .Y(\U1/aes_core/MC3/n98 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U89  ( .A(\U1/aes_core/sb0 [21]), .B(
        \U1/aes_core/sb3 [29]), .Y(\U1/aes_core/MC3/n136 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U88  ( .A(\U1/aes_core/sb2 [5]), .B(
        \U1/aes_core/MC3/n136 ), .Y(\U1/aes_core/MC3/n83 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U87  ( .A(\U1/aes_core/MC3/n98 ), .B(
        \U1/aes_core/MC3/n83 ), .Y(\U1/aes_core/sc3 [13]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U86  ( .A(\U1/aes_core/sb1 [13]), .B(
        \U1/aes_core/sb2 [5]), .Y(\U1/aes_core/MC3/n122 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U85  ( .A(\U1/aes_core/sb0 [22]), .B(
        \U1/aes_core/sb3 [30]), .Y(\U1/aes_core/MC3/n139 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U84  ( .A(\U1/aes_core/sb2 [6]), .B(
        \U1/aes_core/MC3/n139 ), .Y(\U1/aes_core/MC3/n84 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U83  ( .A(\U1/aes_core/MC3/n122 ), .B(
        \U1/aes_core/MC3/n84 ), .Y(\U1/aes_core/sc3 [14]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U82  ( .A(\U1/aes_core/MC3/n142 ), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/MC3/n106 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U81  ( .A(\U1/aes_core/sb1 [14]), .B(
        \U1/aes_core/sb2 [6]), .Y(\U1/aes_core/MC3/n127 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U80  ( .A(\U1/aes_core/sb0 [23]), .B(
        \U1/aes_core/MC3/n127 ), .Y(\U1/aes_core/MC3/n85 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U79  ( .A(\U1/aes_core/MC3/n106 ), .B(
        \U1/aes_core/MC3/n85 ), .Y(\U1/aes_core/sc3 [15]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U78  ( .A(\U1/aes_core/sb3 [24]), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/MC3/n148 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U77  ( .A(\U1/aes_core/sb1 [8]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/MC3/n86 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U76  ( .A(\U1/aes_core/MC3/n86 ), .B(
        \U1/aes_core/sb2 [0]), .Y(\U1/aes_core/MC3/n110 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U75  ( .A(\U1/aes_core/MC3/n148 ), .B(
        \U1/aes_core/MC3/n110 ), .Y(\U1/aes_core/sc3 [16]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U74  ( .A(\U1/aes_core/sb0 [16]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/MC3/n88 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U73  ( .A(\U1/aes_core/MC3/n88 ), .B(
        \U1/aes_core/MC3/n87 ), .Y(\U1/aes_core/MC3/n111 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U72  ( .A(\U1/aes_core/MC3/n89 ), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/MC3/n150 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U71  ( .A(\U1/aes_core/sb3 [25]), .B(
        \U1/aes_core/MC3/n150 ), .Y(\U1/aes_core/MC3/n90 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U70  ( .A(\U1/aes_core/MC3/n111 ), .B(
        \U1/aes_core/MC3/n90 ), .Y(\U1/aes_core/sc3 [17]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U69  ( .A(\U1/aes_core/sb1 [9]), .B(
        \U1/aes_core/sb0 [17]), .Y(\U1/aes_core/MC3/n93 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U68  ( .A(\U1/aes_core/sb1 [10]), .B(
        \U1/aes_core/MC3/n91 ), .Y(\U1/aes_core/MC3/n92 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U67  ( .A(\U1/aes_core/MC3/n93 ), .B(
        \U1/aes_core/MC3/n92 ), .Y(\U1/aes_core/sc3 [18]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U66  ( .A(\U1/aes_core/sb1 [11]), .B(
        \U1/aes_core/sb0 [18]), .Y(\U1/aes_core/MC3/n95 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U65  ( .A(\U1/aes_core/sb2 [3]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/MC3/n94 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U64  ( .A(\U1/aes_core/MC3/n95 ), .B(
        \U1/aes_core/MC3/n94 ), .Y(\U1/aes_core/MC3/n117 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U63  ( .A(\U1/aes_core/MC3/n117 ), .B(
        \U1/aes_core/MC3/n96 ), .Y(\U1/aes_core/sc3 [19]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U62  ( .A(\U1/aes_core/sb3 [24]), .B(
        \U1/aes_core/sb3 [31]), .Y(\U1/aes_core/MC3/n113 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U61  ( .A(\U1/aes_core/sb0 [17]), .B(
        \U1/aes_core/sb3 [25]), .Y(\U1/aes_core/MC3/n114 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U60  ( .A(\U1/aes_core/sb2 [0]), .B(
        \U1/aes_core/sb2 [7]), .Y(\U1/aes_core/MC3/n146 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U59  ( .A(\U1/aes_core/MC3/n114 ), .B(
        \U1/aes_core/MC3/n146 ), .Y(\U1/aes_core/MC3/n149 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U58  ( .A(\U1/aes_core/MC3/n149 ), .B(
        \U1/aes_core/sb1 [9]), .Y(\U1/aes_core/MC3/n97 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U57  ( .A(\U1/aes_core/MC3/n113 ), .B(
        \U1/aes_core/MC3/n97 ), .Y(\U1/aes_core/sc3 [1]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U56  ( .A(\U1/aes_core/sb0 [19]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/MC3/n99 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U55  ( .A(\U1/aes_core/MC3/n99 ), .B(
        \U1/aes_core/MC3/n98 ), .Y(\U1/aes_core/MC3/n118 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U54  ( .A(\U1/aes_core/MC3/n118 ), .B(
        \U1/aes_core/sb3 [28]), .Y(\U1/aes_core/MC3/n100 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U53  ( .A(\U1/aes_core/MC3/n101 ), .B(
        \U1/aes_core/MC3/n100 ), .Y(\U1/aes_core/sc3 [20]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U52  ( .A(\U1/aes_core/sb3 [29]), .B(
        \U1/aes_core/sb0 [20]), .Y(\U1/aes_core/MC3/n103 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U51  ( .A(\U1/aes_core/sb1 [12]), .B(
        \U1/aes_core/MC3/n122 ), .Y(\U1/aes_core/MC3/n102 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U50  ( .A(\U1/aes_core/MC3/n103 ), .B(
        \U1/aes_core/MC3/n102 ), .Y(\U1/aes_core/sc3 [21]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U49  ( .A(\U1/aes_core/sb3 [30]), .B(
        \U1/aes_core/sb0 [21]), .Y(\U1/aes_core/MC3/n105 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U48  ( .A(\U1/aes_core/sb1 [13]), .B(
        \U1/aes_core/MC3/n127 ), .Y(\U1/aes_core/MC3/n104 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U47  ( .A(\U1/aes_core/MC3/n105 ), .B(
        \U1/aes_core/MC3/n104 ), .Y(\U1/aes_core/sc3 [22]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U46  ( .A(\U1/aes_core/sb0 [22]), .B(
        \U1/aes_core/sb1 [15]), .Y(\U1/aes_core/MC3/n108 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U45  ( .A(\U1/aes_core/sb1 [14]), .B(
        \U1/aes_core/MC3/n106 ), .Y(\U1/aes_core/MC3/n107 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U44  ( .A(\U1/aes_core/MC3/n108 ), .B(
        \U1/aes_core/MC3/n107 ), .Y(\U1/aes_core/sc3 [23]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U43  ( .A(\U1/aes_core/MC3/n110 ), .B(
        \U1/aes_core/MC3/n109 ), .Y(\U1/aes_core/sc3 [24]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U42  ( .A(\U1/aes_core/MC3/n111 ), .B(
        \U1/aes_core/sb0 [17]), .Y(\U1/aes_core/MC3/n112 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U41  ( .A(\U1/aes_core/MC3/n113 ), .B(
        \U1/aes_core/MC3/n112 ), .Y(\U1/aes_core/sc3 [25]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U40  ( .A(\U1/aes_core/sb1 [10]), .B(
        \U1/aes_core/sb0 [18]), .Y(\U1/aes_core/MC3/n123 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U39  ( .A(\U1/aes_core/sb2 [2]), .B(
        \U1/aes_core/MC3/n114 ), .Y(\U1/aes_core/MC3/n115 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U38  ( .A(\U1/aes_core/MC3/n123 ), .B(
        \U1/aes_core/MC3/n115 ), .Y(\U1/aes_core/sc3 [26]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U37  ( .A(\U1/aes_core/sb3 [26]), .B(
        \U1/aes_core/sb3 [31]), .Y(\U1/aes_core/MC3/n116 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U36  ( .A(\U1/aes_core/MC3/n116 ), .B(
        \U1/aes_core/sb0 [19]), .Y(\U1/aes_core/MC3/n130 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U32  ( .A(\U1/aes_core/sb3 [27]), .B(
        \U1/aes_core/MC3/n142 ), .Y(\U1/aes_core/MC3/n135 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U31  ( .A(\U1/aes_core/sb0 [20]), .B(
        \U1/aes_core/MC3/n135 ), .Y(\U1/aes_core/MC3/n119 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U29  ( .A(\U1/aes_core/sb0 [21]), .B(
        \U1/aes_core/MC3/n120 ), .Y(\U1/aes_core/MC3/n121 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U28  ( .A(\U1/aes_core/MC3/n122 ), .B(
        \U1/aes_core/MC3/n121 ), .Y(\U1/aes_core/sc3 [29]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U27  ( .A(\U1/aes_core/sb3 [26]), .B(
        \U1/aes_core/sb3 [25]), .Y(\U1/aes_core/MC3/n125 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U26  ( .A(\U1/aes_core/sb2 [1]), .B(
        \U1/aes_core/MC3/n123 ), .Y(\U1/aes_core/MC3/n124 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U25  ( .A(\U1/aes_core/MC3/n125 ), .B(
        \U1/aes_core/MC3/n124 ), .Y(\U1/aes_core/sc3 [2]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U24  ( .A(\U1/aes_core/sb0 [22]), .B(
        \U1/aes_core/MC3/n136 ), .Y(\U1/aes_core/MC3/n126 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U23  ( .A(\U1/aes_core/MC3/n127 ), .B(
        \U1/aes_core/MC3/n126 ), .Y(\U1/aes_core/sc3 [30]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U22  ( .A(\U1/aes_core/sb1 [15]), .B(
        \U1/aes_core/sb0 [23]), .Y(\U1/aes_core/MC3/n143 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U21  ( .A(\U1/aes_core/sb2 [7]), .B(
        \U1/aes_core/MC3/n143 ), .Y(\U1/aes_core/MC3/n128 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U20  ( .A(\U1/aes_core/MC3/n139 ), .B(
        \U1/aes_core/MC3/n128 ), .Y(\U1/aes_core/sc3 [31]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U19  ( .A(\U1/aes_core/sb1 [11]), .B(
        \U1/aes_core/sb3 [27]), .Y(\U1/aes_core/MC3/n132 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U18  ( .A(\U1/aes_core/MC3/n130 ), .B(
        \U1/aes_core/MC3/n129 ), .Y(\U1/aes_core/MC3/n131 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U17  ( .A(\U1/aes_core/MC3/n132 ), .B(
        \U1/aes_core/MC3/n131 ), .Y(\U1/aes_core/sc3 [3]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U16  ( .A(\U1/aes_core/MC3/n133 ), .B(
        \U1/aes_core/sb1 [12]), .Y(\U1/aes_core/MC3/n134 ) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U15  ( .A(\U1/aes_core/MC3/n135 ), .B(
        \U1/aes_core/MC3/n134 ), .Y(\U1/aes_core/sc3 [4]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U14  ( .A(\U1/aes_core/sb2 [4]), .B(
        \U1/aes_core/sb3 [28]), .Y(\U1/aes_core/MC3/n138 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U13  ( .A(\U1/aes_core/sb1 [13]), .B(
        \U1/aes_core/MC3/n136 ), .Y(\U1/aes_core/MC3/n137 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U12  ( .A(\U1/aes_core/MC3/n138 ), .B(
        \U1/aes_core/MC3/n137 ), .Y(\U1/aes_core/sc3 [5]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U11  ( .A(\U1/aes_core/sb2 [5]), .B(
        \U1/aes_core/sb3 [29]), .Y(\U1/aes_core/MC3/n141 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U10  ( .A(\U1/aes_core/sb1 [14]), .B(
        \U1/aes_core/MC3/n139 ), .Y(\U1/aes_core/MC3/n140 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U9  ( .A(\U1/aes_core/MC3/n141 ), .B(
        \U1/aes_core/MC3/n140 ), .Y(\U1/aes_core/sc3 [6]) );
  XNOR2_X0P5M_A12TL \U1/aes_core/MC3/U8  ( .A(\U1/aes_core/sb2 [6]), .B(
        \U1/aes_core/MC3/n142 ), .Y(\U1/aes_core/MC3/n145 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U7  ( .A(\U1/aes_core/sb3 [30]), .B(
        \U1/aes_core/MC3/n143 ), .Y(\U1/aes_core/MC3/n144 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U6  ( .A(\U1/aes_core/MC3/n145 ), .B(
        \U1/aes_core/MC3/n144 ), .Y(\U1/aes_core/sc3 [7]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U5  ( .A(\U1/aes_core/sb0 [16]), .B(
        \U1/aes_core/MC3/n146 ), .Y(\U1/aes_core/MC3/n147 ) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U4  ( .A(\U1/aes_core/MC3/n148 ), .B(
        \U1/aes_core/MC3/n147 ), .Y(\U1/aes_core/sc3 [8]) );
  XOR2_X0P5M_A12TL \U1/aes_core/MC3/U2  ( .A(\U1/aes_core/sb2 [1]), .B(
        \U1/aes_core/MC3/n150 ), .Y(\U1/aes_core/MC3/n151 ) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U136  ( .A(\U1/keyexpantion/ws [0]), .B(
        \U1/rkey [96]), .Y(\U1/rkey_next [96]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U135  ( .A(\U1/rkey_next [96]), .B(
        \U1/rkey [64]), .Y(\U1/rkey_next [64]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U134  ( .A(\U1/rkey_next [64]), .B(
        \U1/rkey [32]), .Y(\U1/rkey_next [32]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U133  ( .A(\U1/rkey [0]), .B(
        \U1/rkey_next [32]), .Y(\U1/rkey_next [0]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U132  ( .A(\U1/keyexpantion/ws [4]), .B(
        \U1/rkey [100]), .Y(\U1/rkey_next [100]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U131  ( .A(\U1/keyexpantion/ws [5]), .B(
        \U1/rkey [101]), .Y(\U1/rkey_next [101]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U130  ( .A(\U1/keyexpantion/ws [6]), .B(
        \U1/rkey [102]), .Y(\U1/rkey_next [102]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U129  ( .A(\U1/keyexpantion/ws [7]), .B(
        \U1/rkey [103]), .Y(\U1/rkey_next [103]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U128  ( .A(\U1/keyexpantion/ws [8]), .B(
        \U1/rkey [104]), .Y(\U1/rkey_next [104]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U127  ( .A(\U1/keyexpantion/ws [9]), .B(
        \U1/rkey [105]), .Y(\U1/rkey_next [105]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U126  ( .A(\U1/keyexpantion/ws [10]), .B(
        \U1/rkey [106]), .Y(\U1/rkey_next [106]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U125  ( .A(\U1/keyexpantion/ws [11]), .B(
        \U1/rkey [107]), .Y(\U1/rkey_next [107]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U124  ( .A(\U1/keyexpantion/ws [12]), .B(
        \U1/rkey [108]), .Y(\U1/rkey_next [108]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U123  ( .A(\U1/keyexpantion/ws [13]), .B(
        \U1/rkey [109]), .Y(\U1/rkey_next [109]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U122  ( .A(\U1/rkey_next [106]), .B(
        \U1/rkey [74]), .Y(\U1/rkey_next [74]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U121  ( .A(\U1/rkey_next [74]), .B(
        \U1/rkey [42]), .Y(\U1/rkey_next [42]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U120  ( .A(\U1/rkey [10]), .B(
        \U1/rkey_next [42]), .Y(\U1/rkey_next [10]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U119  ( .A(\U1/keyexpantion/ws [14]), .B(
        \U1/rkey [110]), .Y(\U1/rkey_next [110]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U118  ( .A(\U1/keyexpantion/ws [15]), .B(
        \U1/rkey [111]), .Y(\U1/rkey_next [111]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U117  ( .A(\U1/keyexpantion/ws [16]), .B(
        \U1/rkey [112]), .Y(\U1/rkey_next [112]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U116  ( .A(\U1/keyexpantion/ws [17]), .B(
        \U1/rkey [113]), .Y(\U1/rkey_next [113]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U115  ( .A(\U1/keyexpantion/ws [18]), .B(
        \U1/rkey [114]), .Y(\U1/rkey_next [114]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U114  ( .A(\U1/keyexpantion/ws [19]), .B(
        \U1/rkey [115]), .Y(\U1/rkey_next [115]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U113  ( .A(\U1/keyexpantion/ws [20]), .B(
        \U1/rkey [116]), .Y(\U1/rkey_next [116]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U112  ( .A(\U1/keyexpantion/ws [21]), .B(
        \U1/rkey [117]), .Y(\U1/rkey_next [117]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U111  ( .A(\U1/keyexpantion/ws [22]), .B(
        \U1/rkey [118]), .Y(\U1/rkey_next [118]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U110  ( .A(\U1/keyexpantion/ws [23]), .B(
        \U1/rkey [119]), .Y(\U1/rkey_next [119]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U109  ( .A(\U1/rkey_next [107]), .B(
        \U1/rkey [75]), .Y(\U1/rkey_next [75]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U108  ( .A(\U1/rkey_next [75]), .B(
        \U1/rkey [43]), .Y(\U1/rkey_next [43]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U107  ( .A(\U1/rkey [11]), .B(
        \U1/rkey_next [43]), .Y(\U1/rkey_next [11]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U106  ( .A(\U1/keyexpantion/ws [24]), .B(
        \U1/rcon [0]), .Y(\U1/keyexpantion/n8 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U105  ( .A(\U1/keyexpantion/n8 ), .B(
        \U1/rkey [120]), .Y(\U1/rkey_next [120]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U104  ( .A(\U1/keyexpantion/ws [25]), .B(
        \U1/rcon [1]), .Y(\U1/keyexpantion/n7 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U103  ( .A(\U1/keyexpantion/n7 ), .B(
        \U1/rkey [121]), .Y(\U1/rkey_next [121]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U102  ( .A(\U1/keyexpantion/ws [26]), .B(
        \U1/rcon [2]), .Y(\U1/keyexpantion/n6 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U101  ( .A(\U1/keyexpantion/n6 ), .B(
        \U1/rkey [122]), .Y(\U1/rkey_next [122]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U100  ( .A(\U1/keyexpantion/ws [27]), .B(
        \U1/rcon [3]), .Y(\U1/keyexpantion/n5 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U99  ( .A(\U1/keyexpantion/n5 ), .B(
        \U1/rkey [123]), .Y(\U1/rkey_next [123]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U98  ( .A(\U1/keyexpantion/ws [28]), .B(
        \U1/rcon [4]), .Y(\U1/keyexpantion/n4 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U97  ( .A(\U1/keyexpantion/n4 ), .B(
        \U1/rkey [124]), .Y(\U1/rkey_next [124]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U96  ( .A(\U1/keyexpantion/ws [29]), .B(
        \U1/rcon [5]), .Y(\U1/keyexpantion/n3 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U95  ( .A(\U1/keyexpantion/n3 ), .B(
        \U1/rkey [125]), .Y(\U1/rkey_next [125]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U94  ( .A(\U1/keyexpantion/ws [30]), .B(
        \U1/rcon [6]), .Y(\U1/keyexpantion/n2 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U93  ( .A(\U1/keyexpantion/n2 ), .B(
        \U1/rkey [126]), .Y(\U1/rkey_next [126]) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U92  ( .A(\U1/keyexpantion/ws [31]), .B(
        \U1/rcon [7]), .Y(\U1/keyexpantion/n1 ) );
  XNOR2_X0P5M_A12TL \U1/keyexpantion/U91  ( .A(\U1/keyexpantion/n1 ), .B(
        \U1/rkey [127]), .Y(\U1/rkey_next [127]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U90  ( .A(\U1/rkey_next [108]), .B(
        \U1/rkey [76]), .Y(\U1/rkey_next [76]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U89  ( .A(\U1/rkey_next [76]), .B(
        \U1/rkey [44]), .Y(\U1/rkey_next [44]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U88  ( .A(\U1/rkey [12]), .B(
        \U1/rkey_next [44]), .Y(\U1/rkey_next [12]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U87  ( .A(\U1/rkey_next [109]), .B(
        \U1/rkey [77]), .Y(\U1/rkey_next [77]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U86  ( .A(\U1/rkey_next [77]), .B(
        \U1/rkey [45]), .Y(\U1/rkey_next [45]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U85  ( .A(\U1/rkey [13]), .B(
        \U1/rkey_next [45]), .Y(\U1/rkey_next [13]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U84  ( .A(\U1/rkey_next [110]), .B(
        \U1/rkey [78]), .Y(\U1/rkey_next [78]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U83  ( .A(\U1/rkey_next [78]), .B(
        \U1/rkey [46]), .Y(\U1/rkey_next [46]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U82  ( .A(\U1/rkey [14]), .B(
        \U1/rkey_next [46]), .Y(\U1/rkey_next [14]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U81  ( .A(\U1/rkey_next [111]), .B(
        \U1/rkey [79]), .Y(\U1/rkey_next [79]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U80  ( .A(\U1/rkey_next [79]), .B(
        \U1/rkey [47]), .Y(\U1/rkey_next [47]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U79  ( .A(\U1/rkey [15]), .B(
        \U1/rkey_next [47]), .Y(\U1/rkey_next [15]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U78  ( .A(\U1/rkey_next [112]), .B(
        \U1/rkey [80]), .Y(\U1/rkey_next [80]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U77  ( .A(\U1/rkey_next [80]), .B(
        \U1/rkey [48]), .Y(\U1/rkey_next [48]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U76  ( .A(\U1/rkey [16]), .B(
        \U1/rkey_next [48]), .Y(\U1/rkey_next [16]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U75  ( .A(\U1/rkey_next [113]), .B(
        \U1/rkey [81]), .Y(\U1/rkey_next [81]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U74  ( .A(\U1/rkey_next [81]), .B(
        \U1/rkey [49]), .Y(\U1/rkey_next [49]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U73  ( .A(\U1/rkey [17]), .B(
        \U1/rkey_next [49]), .Y(\U1/rkey_next [17]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U72  ( .A(\U1/rkey_next [114]), .B(
        \U1/rkey [82]), .Y(\U1/rkey_next [82]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U71  ( .A(\U1/rkey_next [82]), .B(
        \U1/rkey [50]), .Y(\U1/rkey_next [50]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U70  ( .A(\U1/rkey [18]), .B(
        \U1/rkey_next [50]), .Y(\U1/rkey_next [18]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U69  ( .A(\U1/rkey_next [115]), .B(
        \U1/rkey [83]), .Y(\U1/rkey_next [83]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U68  ( .A(\U1/rkey_next [83]), .B(
        \U1/rkey [51]), .Y(\U1/rkey_next [51]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U67  ( .A(\U1/rkey [19]), .B(
        \U1/rkey_next [51]), .Y(\U1/rkey_next [19]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U66  ( .A(\U1/keyexpantion/ws [1]), .B(
        \U1/rkey [97]), .Y(\U1/rkey_next [97]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U65  ( .A(\U1/rkey_next [97]), .B(
        \U1/rkey [65]), .Y(\U1/rkey_next [65]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U64  ( .A(\U1/rkey_next [65]), .B(
        \U1/rkey [33]), .Y(\U1/rkey_next [33]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U63  ( .A(\U1/rkey [1]), .B(
        \U1/rkey_next [33]), .Y(\U1/rkey_next [1]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U62  ( .A(\U1/rkey_next [116]), .B(
        \U1/rkey [84]), .Y(\U1/rkey_next [84]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U61  ( .A(\U1/rkey_next [84]), .B(
        \U1/rkey [52]), .Y(\U1/rkey_next [52]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U60  ( .A(\U1/rkey [20]), .B(
        \U1/rkey_next [52]), .Y(\U1/rkey_next [20]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U59  ( .A(\U1/rkey_next [117]), .B(
        \U1/rkey [85]), .Y(\U1/rkey_next [85]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U58  ( .A(\U1/rkey_next [85]), .B(
        \U1/rkey [53]), .Y(\U1/rkey_next [53]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U57  ( .A(\U1/rkey [21]), .B(
        \U1/rkey_next [53]), .Y(\U1/rkey_next [21]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U56  ( .A(\U1/rkey_next [118]), .B(
        \U1/rkey [86]), .Y(\U1/rkey_next [86]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U55  ( .A(\U1/rkey_next [86]), .B(
        \U1/rkey [54]), .Y(\U1/rkey_next [54]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U54  ( .A(\U1/rkey [22]), .B(
        \U1/rkey_next [54]), .Y(\U1/rkey_next [22]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U53  ( .A(\U1/rkey_next [119]), .B(
        \U1/rkey [87]), .Y(\U1/rkey_next [87]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U52  ( .A(\U1/rkey_next [87]), .B(
        \U1/rkey [55]), .Y(\U1/rkey_next [55]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U51  ( .A(\U1/rkey [23]), .B(
        \U1/rkey_next [55]), .Y(\U1/rkey_next [23]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U50  ( .A(\U1/rkey_next [120]), .B(
        \U1/rkey [88]), .Y(\U1/rkey_next [88]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U49  ( .A(\U1/rkey_next [88]), .B(
        \U1/rkey [56]), .Y(\U1/rkey_next [56]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U48  ( .A(\U1/rkey [24]), .B(
        \U1/rkey_next [56]), .Y(\U1/rkey_next [24]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U47  ( .A(\U1/rkey_next [121]), .B(
        \U1/rkey [89]), .Y(\U1/rkey_next [89]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U46  ( .A(\U1/rkey_next [89]), .B(
        \U1/rkey [57]), .Y(\U1/rkey_next [57]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U45  ( .A(\U1/rkey [25]), .B(
        \U1/rkey_next [57]), .Y(\U1/rkey_next [25]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U44  ( .A(\U1/rkey_next [122]), .B(
        \U1/rkey [90]), .Y(\U1/rkey_next [90]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U43  ( .A(\U1/rkey_next [90]), .B(
        \U1/rkey [58]), .Y(\U1/rkey_next [58]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U42  ( .A(\U1/rkey [26]), .B(
        \U1/rkey_next [58]), .Y(\U1/rkey_next [26]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U41  ( .A(\U1/rkey_next [123]), .B(
        \U1/rkey [91]), .Y(\U1/rkey_next [91]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U40  ( .A(\U1/rkey_next [91]), .B(
        \U1/rkey [59]), .Y(\U1/rkey_next [59]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U39  ( .A(\U1/rkey [27]), .B(
        \U1/rkey_next [59]), .Y(\U1/rkey_next [27]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U38  ( .A(\U1/rkey_next [124]), .B(
        \U1/rkey [92]), .Y(\U1/rkey_next [92]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U37  ( .A(\U1/rkey_next [92]), .B(
        \U1/rkey [60]), .Y(\U1/rkey_next [60]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U36  ( .A(\U1/rkey [28]), .B(
        \U1/rkey_next [60]), .Y(\U1/rkey_next [28]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U35  ( .A(\U1/rkey_next [125]), .B(
        \U1/rkey [93]), .Y(\U1/rkey_next [93]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U34  ( .A(\U1/rkey_next [93]), .B(
        \U1/rkey [61]), .Y(\U1/rkey_next [61]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U33  ( .A(\U1/rkey [29]), .B(
        \U1/rkey_next [61]), .Y(\U1/rkey_next [29]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U32  ( .A(\U1/keyexpantion/ws [2]), .B(
        \U1/rkey [98]), .Y(\U1/rkey_next [98]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U31  ( .A(\U1/rkey_next [98]), .B(
        \U1/rkey [66]), .Y(\U1/rkey_next [66]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U30  ( .A(\U1/rkey_next [66]), .B(
        \U1/rkey [34]), .Y(\U1/rkey_next [34]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U29  ( .A(\U1/rkey [2]), .B(
        \U1/rkey_next [34]), .Y(\U1/rkey_next [2]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U28  ( .A(\U1/rkey_next [126]), .B(
        \U1/rkey [94]), .Y(\U1/rkey_next [94]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U27  ( .A(\U1/rkey_next [94]), .B(
        \U1/rkey [62]), .Y(\U1/rkey_next [62]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U26  ( .A(\U1/rkey [30]), .B(
        \U1/rkey_next [62]), .Y(\U1/rkey_next [30]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U25  ( .A(\U1/rkey_next [127]), .B(
        \U1/rkey [95]), .Y(\U1/rkey_next [95]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U24  ( .A(\U1/rkey_next [95]), .B(
        \U1/rkey [63]), .Y(\U1/rkey_next [63]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U23  ( .A(\U1/rkey [31]), .B(
        \U1/rkey_next [63]), .Y(\U1/rkey_next [31]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U22  ( .A(\U1/keyexpantion/ws [3]), .B(
        \U1/rkey [99]), .Y(\U1/rkey_next [99]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U21  ( .A(\U1/rkey_next [99]), .B(
        \U1/rkey [67]), .Y(\U1/rkey_next [67]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U20  ( .A(\U1/rkey_next [67]), .B(
        \U1/rkey [35]), .Y(\U1/rkey_next [35]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U19  ( .A(\U1/rkey_next [100]), .B(
        \U1/rkey [68]), .Y(\U1/rkey_next [68]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U18  ( .A(\U1/rkey_next [68]), .B(
        \U1/rkey [36]), .Y(\U1/rkey_next [36]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U17  ( .A(\U1/rkey_next [101]), .B(
        \U1/rkey [69]), .Y(\U1/rkey_next [69]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U16  ( .A(\U1/rkey_next [69]), .B(
        \U1/rkey [37]), .Y(\U1/rkey_next [37]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U15  ( .A(\U1/rkey_next [102]), .B(
        \U1/rkey [70]), .Y(\U1/rkey_next [70]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U14  ( .A(\U1/rkey_next [70]), .B(
        \U1/rkey [38]), .Y(\U1/rkey_next [38]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U13  ( .A(\U1/rkey_next [103]), .B(
        \U1/rkey [71]), .Y(\U1/rkey_next [71]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U12  ( .A(\U1/rkey_next [71]), .B(
        \U1/rkey [39]), .Y(\U1/rkey_next [39]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U11  ( .A(\U1/rkey [3]), .B(
        \U1/rkey_next [35]), .Y(\U1/rkey_next [3]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U10  ( .A(\U1/rkey_next [104]), .B(
        \U1/rkey [72]), .Y(\U1/rkey_next [72]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U9  ( .A(\U1/rkey_next [72]), .B(
        \U1/rkey [40]), .Y(\U1/rkey_next [40]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U8  ( .A(\U1/rkey_next [105]), .B(
        \U1/rkey [73]), .Y(\U1/rkey_next [73]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U7  ( .A(\U1/rkey_next [73]), .B(
        \U1/rkey [41]), .Y(\U1/rkey_next [41]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U6  ( .A(\U1/rkey [4]), .B(
        \U1/rkey_next [36]), .Y(\U1/rkey_next [4]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U5  ( .A(\U1/rkey [5]), .B(
        \U1/rkey_next [37]), .Y(\U1/rkey_next [5]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U4  ( .A(\U1/rkey [6]), .B(
        \U1/rkey_next [38]), .Y(\U1/rkey_next [6]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U3  ( .A(\U1/rkey [7]), .B(
        \U1/rkey_next [39]), .Y(\U1/rkey_next [7]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U2  ( .A(\U1/rkey [8]), .B(
        \U1/rkey_next [40]), .Y(\U1/rkey_next [8]) );
  XOR2_X0P5M_A12TL \U1/keyexpantion/U1  ( .A(\U1/rkey [9]), .B(
        \U1/rkey_next [41]), .Y(\U1/rkey_next [9]) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U363  ( .A0(
        \U1/keyexpantion/SB0/n2833 ), .A1(\U1/keyexpantion/SB0/n2613 ), .B0(
        \U1/keyexpantion/SB0/n2932 ), .B1(\U1/keyexpantion/SB0/n2916 ), .C0(
        \U1/keyexpantion/SB0/n2681 ), .Y(\U1/keyexpantion/SB0/n2614 ) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U361  ( .A0(
        \U1/keyexpantion/SB0/n2211 ), .A1(\U1/keyexpantion/SB0/n2361 ), .B0(
        \U1/keyexpantion/SB0/n2359 ), .B1(\U1/keyexpantion/SB0/n2319 ), .C0(
        \U1/keyexpantion/SB0/n2210 ), .Y(\U1/keyexpantion/SB0/n2213 ) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U301  ( .A0(
        \U1/keyexpantion/SB0/n2980 ), .A1(\U1/keyexpantion/SB0/n3105 ), .B0(
        \U1/keyexpantion/SB0/n3103 ), .B1(\U1/keyexpantion/SB0/n3088 ), .C0(
        \U1/keyexpantion/SB0/n2979 ), .Y(\U1/keyexpantion/SB0/n2982 ) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U300  ( .A0(
        \U1/keyexpantion/SB0/n2410 ), .A1(\U1/keyexpantion/SB0/n2165 ), .B0(
        \U1/keyexpantion/SB0/n2488 ), .B1(\U1/keyexpantion/SB0/n2472 ), .C0(
        \U1/keyexpantion/SB0/n2233 ), .Y(\U1/keyexpantion/SB0/n2166 ) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U151  ( .A0(
        \U1/keyexpantion/SB0/n3154 ), .A1(\U1/keyexpantion/SB0/n2336 ), .B0(
        \U1/keyexpantion/SB0/n3232 ), .B1(\U1/keyexpantion/SB0/n3216 ), .C0(
        \U1/keyexpantion/SB0/n3002 ), .Y(\U1/keyexpantion/SB0/n2337 ) );
  OAI221_X1M_A12TL \U1/keyexpantion/SB0/U150  ( .A0(
        \U1/keyexpantion/SB0/n2659 ), .A1(\U1/keyexpantion/SB0/n2784 ), .B0(
        \U1/keyexpantion/SB0/n2782 ), .B1(\U1/keyexpantion/SB0/n2767 ), .C0(
        \U1/keyexpantion/SB0/n2658 ), .Y(\U1/keyexpantion/SB0/n2661 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1724  ( .A(\U1/rkey [31]), .B(
        \U1/rkey [30]), .Y(\U1/keyexpantion/SB0/n1697 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1723  ( .A(\U1/rkey [29]), .B(
        \U1/rkey [28]), .Y(\U1/keyexpantion/SB0/n1688 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1722  ( .A(
        \U1/keyexpantion/SB0/n1697 ), .B(\U1/keyexpantion/SB0/n1688 ), .Y(
        \U1/keyexpantion/SB0/n2336 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1721  ( .A(\U1/rkey [25]), .Y(
        \U1/keyexpantion/SB0/n1030 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1720  ( .A(\U1/rkey [24]), .Y(
        \U1/keyexpantion/SB0/n385 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1719  ( .A(
        \U1/keyexpantion/SB0/n1030 ), .B(\U1/keyexpantion/SB0/n385 ), .Y(
        \U1/keyexpantion/SB0/n1689 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1718  ( .A(\U1/rkey [27]), .B(
        \U1/rkey [26]), .Y(\U1/keyexpantion/SB0/n1709 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1717  ( .A(
        \U1/keyexpantion/SB0/n1689 ), .B(\U1/keyexpantion/SB0/n1709 ), .Y(
        \U1/keyexpantion/SB0/n3216 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1716  ( .A(
        \U1/keyexpantion/SB0/n2336 ), .B(\U1/keyexpantion/SB0/n3216 ), .Y(
        \U1/keyexpantion/SB0/n3023 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U1715  ( .A(\U1/rkey [26]), .B(
        \U1/rkey [27]), .Y(\U1/keyexpantion/SB0/n1692 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1714  ( .A(
        \U1/keyexpantion/SB0/n1692 ), .B(\U1/keyexpantion/SB0/n1689 ), .Y(
        \U1/keyexpantion/SB0/n3154 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1713  ( .A(\U1/rkey [31]), .Y(
        \U1/keyexpantion/SB0/n1685 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1712  ( .A(
        \U1/keyexpantion/SB0/n1685 ), .B(\U1/rkey [30]), .Y(
        \U1/keyexpantion/SB0/n1715 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1711  ( .A(
        \U1/keyexpantion/SB0/n1715 ), .B(\U1/keyexpantion/SB0/n1688 ), .Y(
        \U1/keyexpantion/SB0/n2335 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1710  ( .A(
        \U1/keyexpantion/SB0/n3154 ), .B(\U1/keyexpantion/SB0/n2335 ), .Y(
        \U1/keyexpantion/SB0/n3120 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1709  ( .A(\U1/rkey [27]), .Y(
        \U1/keyexpantion/SB0/n707 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U1708  ( .A(\U1/rkey [26]), .B(
        \U1/keyexpantion/SB0/n707 ), .Y(\U1/keyexpantion/SB0/n1690 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1707  ( .A(
        \U1/keyexpantion/SB0/n1689 ), .B(\U1/keyexpantion/SB0/n1690 ), .Y(
        \U1/keyexpantion/SB0/n3085 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1706  ( .A(\U1/keyexpantion/SB0/n3085 ), .Y(\U1/keyexpantion/SB0/n3250 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1705  ( .A(\U1/rkey [28]), .Y(
        \U1/keyexpantion/SB0/n752 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1704  ( .A(\U1/keyexpantion/SB0/n752 ), .B(\U1/rkey [29]), .Y(\U1/keyexpantion/SB0/n1696 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1703  ( .A(\U1/rkey [30]), .Y(
        \U1/keyexpantion/SB0/n1203 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1702  ( .A(
        \U1/keyexpantion/SB0/n1203 ), .B(\U1/rkey [31]), .Y(
        \U1/keyexpantion/SB0/n1706 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1701  ( .A(
        \U1/keyexpantion/SB0/n1696 ), .B(\U1/keyexpantion/SB0/n1706 ), .Y(
        \U1/keyexpantion/SB0/n3106 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1700  ( .A(\U1/keyexpantion/SB0/n3106 ), .Y(\U1/keyexpantion/SB0/n3204 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1699  ( .A(
        \U1/keyexpantion/SB0/n3250 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3063 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1698  ( .A(\U1/keyexpantion/SB0/n2336 ), .Y(\U1/keyexpantion/SB0/n3219 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1697  ( .A(\U1/rkey [25]), .B(
        \U1/rkey [24]), .Y(\U1/keyexpantion/SB0/n1693 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1696  ( .A(
        \U1/keyexpantion/SB0/n1693 ), .B(\U1/keyexpantion/SB0/n1709 ), .Y(
        \U1/keyexpantion/SB0/n3172 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1695  ( .A(\U1/keyexpantion/SB0/n3172 ), .Y(\U1/keyexpantion/SB0/n3260 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1694  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3260 ), .Y(
        \U1/keyexpantion/SB0/n3177 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1693  ( .A(\U1/keyexpantion/SB0/n385 ), .B(\U1/rkey [25]), .Y(\U1/keyexpantion/SB0/n1708 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1692  ( .A(
        \U1/keyexpantion/SB0/n1690 ), .B(\U1/keyexpantion/SB0/n1708 ), .Y(
        \U1/keyexpantion/SB0/n3072 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1691  ( .A(\U1/keyexpantion/SB0/n3072 ), .Y(\U1/keyexpantion/SB0/n3161 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1690  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3041 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U1689  ( .A(
        \U1/keyexpantion/SB0/n3063 ), .B(\U1/keyexpantion/SB0/n3177 ), .C(
        \U1/keyexpantion/SB0/n3041 ), .Y(\U1/keyexpantion/SB0/n1728 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1688  ( .A(
        \U1/keyexpantion/SB0/n1688 ), .B(\U1/keyexpantion/SB0/n1706 ), .Y(
        \U1/keyexpantion/SB0/n3105 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1687  ( .A(\U1/keyexpantion/SB0/n707 ), .B(\U1/rkey [26]), .Y(\U1/keyexpantion/SB0/n1699 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1686  ( .A(
        \U1/keyexpantion/SB0/n1699 ), .B(\U1/keyexpantion/SB0/n1708 ), .Y(
        \U1/keyexpantion/SB0/n3103 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1685  ( .A(
        \U1/keyexpantion/SB0/n3105 ), .B(\U1/keyexpantion/SB0/n3103 ), .Y(
        \U1/keyexpantion/SB0/n3018 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1684  ( .A(\U1/keyexpantion/SB0/n2335 ), .Y(\U1/keyexpantion/SB0/n3221 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1683  ( .A(\U1/rkey [29]), .Y(
        \U1/keyexpantion/SB0/n1158 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1682  ( .A(\U1/keyexpantion/SB0/n752 ), .B(\U1/keyexpantion/SB0/n1158 ), .Y(\U1/keyexpantion/SB0/n1707 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1681  ( .A(
        \U1/keyexpantion/SB0/n1697 ), .B(\U1/keyexpantion/SB0/n1707 ), .Y(
        \U1/keyexpantion/SB0/n3264 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1680  ( .A(\U1/keyexpantion/SB0/n3264 ), .Y(\U1/keyexpantion/SB0/n3195 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1679  ( .A(
        \U1/keyexpantion/SB0/n1030 ), .B(\U1/rkey [24]), .Y(
        \U1/keyexpantion/SB0/n1698 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1678  ( .A(
        \U1/keyexpantion/SB0/n1698 ), .B(\U1/keyexpantion/SB0/n1709 ), .Y(
        \U1/keyexpantion/SB0/n3229 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1677  ( .A(\U1/keyexpantion/SB0/n3229 ), .Y(\U1/keyexpantion/SB0/n3077 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1676  ( .A0(
        \U1/keyexpantion/SB0/n3221 ), .A1(\U1/keyexpantion/SB0/n3195 ), .B0(
        \U1/keyexpantion/SB0/n3077 ), .Y(\U1/keyexpantion/SB0/n1687 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1675  ( .A(
        \U1/keyexpantion/SB0/n1693 ), .B(\U1/keyexpantion/SB0/n1690 ), .Y(
        \U1/keyexpantion/SB0/n3217 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1674  ( .A(\U1/keyexpantion/SB0/n3217 ), .Y(\U1/keyexpantion/SB0/n3203 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1673  ( .A(
        \U1/keyexpantion/SB0/n1158 ), .B(\U1/rkey [28]), .Y(
        \U1/keyexpantion/SB0/n1714 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1672  ( .A(
        \U1/keyexpantion/SB0/n1706 ), .B(\U1/keyexpantion/SB0/n1714 ), .Y(
        \U1/keyexpantion/SB0/n3257 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1671  ( .A(
        \U1/keyexpantion/SB0/n3105 ), .B(\U1/keyexpantion/SB0/n3257 ), .Y(
        \U1/keyexpantion/SB0/n2996 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1670  ( .A(
        \U1/keyexpantion/SB0/n1685 ), .B(\U1/keyexpantion/SB0/n1203 ), .Y(
        \U1/keyexpantion/SB0/n1705 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1669  ( .A(
        \U1/keyexpantion/SB0/n1696 ), .B(\U1/keyexpantion/SB0/n1705 ), .Y(
        \U1/keyexpantion/SB0/n3232 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1668  ( .A(\U1/keyexpantion/SB0/n3232 ), .Y(\U1/keyexpantion/SB0/n2977 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1667  ( .A0(
        \U1/keyexpantion/SB0/n3203 ), .A1(\U1/keyexpantion/SB0/n2996 ), .B0(
        \U1/keyexpantion/SB0/n2977 ), .B1(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n1686 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1666  ( .AN(
        \U1/keyexpantion/SB0/n3018 ), .B(\U1/keyexpantion/SB0/n1687 ), .C(
        \U1/keyexpantion/SB0/n1686 ), .Y(\U1/keyexpantion/SB0/n1727 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1665  ( .A(
        \U1/keyexpantion/SB0/n1688 ), .B(\U1/keyexpantion/SB0/n1705 ), .Y(
        \U1/keyexpantion/SB0/n3122 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1664  ( .A(
        \U1/keyexpantion/SB0/n1692 ), .B(\U1/keyexpantion/SB0/n1693 ), .Y(
        \U1/keyexpantion/SB0/n3267 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1663  ( .A(
        \U1/keyexpantion/SB0/n1715 ), .B(\U1/keyexpantion/SB0/n1696 ), .Y(
        \U1/keyexpantion/SB0/n3173 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1662  ( .A(
        \U1/keyexpantion/SB0/n1692 ), .B(\U1/keyexpantion/SB0/n1698 ), .Y(
        \U1/keyexpantion/SB0/n3170 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1661  ( .A(
        \U1/keyexpantion/SB0/n1689 ), .B(\U1/keyexpantion/SB0/n1699 ), .Y(
        \U1/keyexpantion/SB0/n3175 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1660  ( .A(\U1/keyexpantion/SB0/n3175 ), .Y(\U1/keyexpantion/SB0/n3155 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1659  ( .A(\U1/keyexpantion/SB0/n3257 ), .Y(\U1/keyexpantion/SB0/n2991 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1658  ( .A(
        \U1/keyexpantion/SB0/n1690 ), .B(\U1/keyexpantion/SB0/n1698 ), .Y(
        \U1/keyexpantion/SB0/n3193 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1657  ( .A(\U1/keyexpantion/SB0/n3193 ), .Y(\U1/keyexpantion/SB0/n3218 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1656  ( .A0(
        \U1/keyexpantion/SB0/n3155 ), .A1(\U1/keyexpantion/SB0/n3219 ), .B0(
        \U1/keyexpantion/SB0/n2991 ), .B1(\U1/keyexpantion/SB0/n3218 ), .Y(
        \U1/keyexpantion/SB0/n1691 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1655  ( .A0(
        \U1/keyexpantion/SB0/n3122 ), .A1(\U1/keyexpantion/SB0/n3267 ), .B0(
        \U1/keyexpantion/SB0/n3173 ), .B1(\U1/keyexpantion/SB0/n3170 ), .C0(
        \U1/keyexpantion/SB0/n1691 ), .Y(\U1/keyexpantion/SB0/n1726 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1654  ( .A(
        \U1/keyexpantion/SB0/n3175 ), .B(\U1/keyexpantion/SB0/n3122 ), .Y(
        \U1/keyexpantion/SB0/n2984 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1653  ( .A(
        \U1/keyexpantion/SB0/n3170 ), .B(\U1/keyexpantion/SB0/n3105 ), .Y(
        \U1/keyexpantion/SB0/n2994 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1652  ( .A(\U1/keyexpantion/SB0/n2994 ), .Y(\U1/keyexpantion/SB0/n1695 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1651  ( .A(
        \U1/keyexpantion/SB0/n1692 ), .B(\U1/keyexpantion/SB0/n1708 ), .Y(
        \U1/keyexpantion/SB0/n3245 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1650  ( .A(\U1/keyexpantion/SB0/n3245 ), .Y(\U1/keyexpantion/SB0/n3194 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1649  ( .A(
        \U1/keyexpantion/SB0/n1693 ), .B(\U1/keyexpantion/SB0/n1699 ), .Y(
        \U1/keyexpantion/SB0/n3230 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1648  ( .A(\U1/keyexpantion/SB0/n3230 ), .Y(\U1/keyexpantion/SB0/n3241 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1647  ( .A0(
        \U1/keyexpantion/SB0/n3194 ), .A1(\U1/keyexpantion/SB0/n3241 ), .B0(
        \U1/keyexpantion/SB0/n3195 ), .Y(\U1/keyexpantion/SB0/n1694 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1646  ( .A(
        \U1/keyexpantion/SB0/n1697 ), .B(\U1/keyexpantion/SB0/n1714 ), .Y(
        \U1/keyexpantion/SB0/n3246 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1645  ( .A(\U1/keyexpantion/SB0/n3246 ), .Y(\U1/keyexpantion/SB0/n3196 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1644  ( .A(
        \U1/keyexpantion/SB0/n3196 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3011 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1643  ( .AN(
        \U1/keyexpantion/SB0/n2984 ), .B(\U1/keyexpantion/SB0/n1695 ), .C(
        \U1/keyexpantion/SB0/n1694 ), .D(\U1/keyexpantion/SB0/n3011 ), .Y(
        \U1/keyexpantion/SB0/n1704 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1642  ( .A(
        \U1/keyexpantion/SB0/n1707 ), .B(\U1/keyexpantion/SB0/n1705 ), .Y(
        \U1/keyexpantion/SB0/n3266 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1641  ( .A(
        \U1/keyexpantion/SB0/n1697 ), .B(\U1/keyexpantion/SB0/n1696 ), .Y(
        \U1/keyexpantion/SB0/n3258 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1640  ( .A0(
        \U1/keyexpantion/SB0/n2335 ), .A1(\U1/keyexpantion/SB0/n3085 ), .B0(
        \U1/keyexpantion/SB0/n3266 ), .B1(\U1/keyexpantion/SB0/n3175 ), .C0(
        \U1/keyexpantion/SB0/n3258 ), .C1(\U1/keyexpantion/SB0/n3193 ), .Y(
        \U1/keyexpantion/SB0/n1703 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1639  ( .A(
        \U1/keyexpantion/SB0/n3217 ), .B(\U1/keyexpantion/SB0/n2335 ), .Y(
        \U1/keyexpantion/SB0/n3069 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1638  ( .A(
        \U1/keyexpantion/SB0/n2991 ), .B(\U1/keyexpantion/SB0/n3155 ), .Y(
        \U1/keyexpantion/SB0/n3022 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1637  ( .A(
        \U1/keyexpantion/SB0/n3218 ), .B(\U1/keyexpantion/SB0/n3219 ), .Y(
        \U1/keyexpantion/SB0/n3042 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1636  ( .A(\U1/keyexpantion/SB0/n3173 ), .Y(\U1/keyexpantion/SB0/n3247 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1635  ( .A(
        \U1/keyexpantion/SB0/n3247 ), .B(\U1/keyexpantion/SB0/n3077 ), .Y(
        \U1/keyexpantion/SB0/n3080 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1634  ( .AN(
        \U1/keyexpantion/SB0/n3069 ), .B(\U1/keyexpantion/SB0/n3022 ), .C(
        \U1/keyexpantion/SB0/n3042 ), .D(\U1/keyexpantion/SB0/n3080 ), .Y(
        \U1/keyexpantion/SB0/n1702 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1633  ( .A(
        \U1/keyexpantion/SB0/n1715 ), .B(\U1/keyexpantion/SB0/n1707 ), .Y(
        \U1/keyexpantion/SB0/n2992 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1632  ( .A(
        \U1/keyexpantion/SB0/n2992 ), .B(\U1/keyexpantion/SB0/n3229 ), .Y(
        \U1/keyexpantion/SB0/n3146 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1631  ( .A(
        \U1/keyexpantion/SB0/n1699 ), .B(\U1/keyexpantion/SB0/n1698 ), .Y(
        \U1/keyexpantion/SB0/n3265 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1630  ( .A(
        \U1/keyexpantion/SB0/n3232 ), .B(\U1/keyexpantion/SB0/n3265 ), .Y(
        \U1/keyexpantion/SB0/n3111 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1629  ( .A(\U1/keyexpantion/SB0/n3111 ), .Y(\U1/keyexpantion/SB0/n1700 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1628  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3077 ), .Y(
        \U1/keyexpantion/SB0/n3130 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1627  ( .A(\U1/keyexpantion/SB0/n3265 ), .Y(\U1/keyexpantion/SB0/n3248 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1626  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3248 ), .Y(
        \U1/keyexpantion/SB0/n3181 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1625  ( .AN(
        \U1/keyexpantion/SB0/n3146 ), .B(\U1/keyexpantion/SB0/n1700 ), .C(
        \U1/keyexpantion/SB0/n3130 ), .D(\U1/keyexpantion/SB0/n3181 ), .Y(
        \U1/keyexpantion/SB0/n1701 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1624  ( .A(\U1/keyexpantion/SB0/n1704 ), .B(\U1/keyexpantion/SB0/n1703 ), .C(\U1/keyexpantion/SB0/n1702 ), .D(
        \U1/keyexpantion/SB0/n1701 ), .Y(\U1/keyexpantion/SB0/n2914 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1623  ( .A(
        \U1/keyexpantion/SB0/n3172 ), .B(\U1/keyexpantion/SB0/n2992 ), .Y(
        \U1/keyexpantion/SB0/n3180 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1622  ( .A(
        \U1/keyexpantion/SB0/n1714 ), .B(\U1/keyexpantion/SB0/n1705 ), .Y(
        \U1/keyexpantion/SB0/n3088 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1621  ( .A(
        \U1/keyexpantion/SB0/n3154 ), .B(\U1/keyexpantion/SB0/n3088 ), .Y(
        \U1/keyexpantion/SB0/n3059 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1620  ( .A(\U1/keyexpantion/SB0/n3266 ), .Y(\U1/keyexpantion/SB0/n3222 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1619  ( .A(
        \U1/keyexpantion/SB0/n3222 ), .B(\U1/keyexpantion/SB0/n3203 ), .Y(
        \U1/keyexpantion/SB0/n3008 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1618  ( .A0(
        \U1/keyexpantion/SB0/n3088 ), .A1(\U1/keyexpantion/SB0/n3265 ), .B0(
        \U1/keyexpantion/SB0/n3008 ), .Y(\U1/keyexpantion/SB0/n1713 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1617  ( .A(\U1/keyexpantion/SB0/n3103 ), .Y(\U1/keyexpantion/SB0/n3198 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1616  ( .A(
        \U1/keyexpantion/SB0/n3198 ), .B(\U1/keyexpantion/SB0/n3221 ), .Y(
        \U1/keyexpantion/SB0/n3199 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1615  ( .A(
        \U1/keyexpantion/SB0/n3221 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3158 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1614  ( .A(
        \U1/keyexpantion/SB0/n1707 ), .B(\U1/keyexpantion/SB0/n1706 ), .Y(
        \U1/keyexpantion/SB0/n3228 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1613  ( .A(\U1/keyexpantion/SB0/n3228 ), .Y(\U1/keyexpantion/SB0/n3003 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1612  ( .A(
        \U1/keyexpantion/SB0/n3194 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3027 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1611  ( .A(\U1/keyexpantion/SB0/n3216 ), .Y(\U1/keyexpantion/SB0/n3197 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1610  ( .A(
        \U1/keyexpantion/SB0/n3197 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3091 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1609  ( .A(
        \U1/keyexpantion/SB0/n3199 ), .B(\U1/keyexpantion/SB0/n3158 ), .C(
        \U1/keyexpantion/SB0/n3027 ), .D(\U1/keyexpantion/SB0/n3091 ), .Y(
        \U1/keyexpantion/SB0/n1712 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1608  ( .A(
        \U1/keyexpantion/SB0/n3218 ), .B(\U1/keyexpantion/SB0/n3196 ), .Y(
        \U1/keyexpantion/SB0/n3125 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1607  ( .A(
        \U1/keyexpantion/SB0/n3260 ), .B(\U1/keyexpantion/SB0/n3196 ), .Y(
        \U1/keyexpantion/SB0/n3116 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1606  ( .A(\U1/keyexpantion/SB0/n3258 ), .Y(\U1/keyexpantion/SB0/n3251 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1605  ( .A(
        \U1/keyexpantion/SB0/n3155 ), .B(\U1/keyexpantion/SB0/n3251 ), .Y(
        \U1/keyexpantion/SB0/n2988 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1604  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3194 ), .Y(
        \U1/keyexpantion/SB0/n3099 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1603  ( .A(
        \U1/keyexpantion/SB0/n3125 ), .B(\U1/keyexpantion/SB0/n3116 ), .C(
        \U1/keyexpantion/SB0/n2988 ), .D(\U1/keyexpantion/SB0/n3099 ), .Y(
        \U1/keyexpantion/SB0/n1711 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1602  ( .A(\U1/keyexpantion/SB0/n3170 ), .Y(\U1/keyexpantion/SB0/n3139 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1601  ( .A(
        \U1/keyexpantion/SB0/n2991 ), .B(\U1/keyexpantion/SB0/n3139 ), .Y(
        \U1/keyexpantion/SB0/n2975 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1600  ( .A(
        \U1/keyexpantion/SB0/n1709 ), .B(\U1/keyexpantion/SB0/n1708 ), .Y(
        \U1/keyexpantion/SB0/n3205 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1599  ( .A(\U1/keyexpantion/SB0/n3205 ), .Y(\U1/keyexpantion/SB0/n3239 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1598  ( .A(
        \U1/keyexpantion/SB0/n2991 ), .B(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3039 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1597  ( .A(\U1/keyexpantion/SB0/n3154 ), .Y(\U1/keyexpantion/SB0/n3262 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1596  ( .A(
        \U1/keyexpantion/SB0/n3262 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3074 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1595  ( .A(
        \U1/keyexpantion/SB0/n3195 ), .B(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3223 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1594  ( .A(
        \U1/keyexpantion/SB0/n2975 ), .B(\U1/keyexpantion/SB0/n3039 ), .C(
        \U1/keyexpantion/SB0/n3074 ), .D(\U1/keyexpantion/SB0/n3223 ), .Y(
        \U1/keyexpantion/SB0/n1710 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1593  ( .A(\U1/keyexpantion/SB0/n3180 ), .B(\U1/keyexpantion/SB0/n3059 ), .C(\U1/keyexpantion/SB0/n1713 ), .D(
        \U1/keyexpantion/SB0/n1712 ), .E(\U1/keyexpantion/SB0/n1711 ), .F(
        \U1/keyexpantion/SB0/n1710 ), .Y(\U1/keyexpantion/SB0/n2903 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1592  ( .A(\U1/keyexpantion/SB0/n2903 ), .Y(\U1/keyexpantion/SB0/n1724 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1591  ( .A(
        \U1/keyexpantion/SB0/n3230 ), .B(\U1/keyexpantion/SB0/n3088 ), .Y(
        \U1/keyexpantion/SB0/n2985 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1590  ( .A(
        \U1/keyexpantion/SB0/n1715 ), .B(\U1/keyexpantion/SB0/n1714 ), .Y(
        \U1/keyexpantion/SB0/n3227 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1589  ( .A(
        \U1/keyexpantion/SB0/n3227 ), .B(\U1/keyexpantion/SB0/n3103 ), .Y(
        \U1/keyexpantion/SB0/n3112 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1588  ( .A(\U1/keyexpantion/SB0/n3112 ), .Y(\U1/keyexpantion/SB0/n1717 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1587  ( .A(\U1/keyexpantion/SB0/n3105 ), .Y(\U1/keyexpantion/SB0/n3252 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1586  ( .A0(
        \U1/keyexpantion/SB0/n3003 ), .A1(\U1/keyexpantion/SB0/n3252 ), .B0(
        \U1/keyexpantion/SB0/n3239 ), .Y(\U1/keyexpantion/SB0/n1716 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1585  ( .A(
        \U1/keyexpantion/SB0/n3222 ), .B(\U1/keyexpantion/SB0/n3139 ), .Y(
        \U1/keyexpantion/SB0/n3010 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1584  ( .AN(
        \U1/keyexpantion/SB0/n2985 ), .B(\U1/keyexpantion/SB0/n1717 ), .C(
        \U1/keyexpantion/SB0/n1716 ), .D(\U1/keyexpantion/SB0/n3010 ), .Y(
        \U1/keyexpantion/SB0/n1721 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1583  ( .A0(
        \U1/keyexpantion/SB0/n3216 ), .A1(\U1/keyexpantion/SB0/n3264 ), .B0(
        \U1/keyexpantion/SB0/n3122 ), .B1(\U1/keyexpantion/SB0/n3170 ), .C0(
        \U1/keyexpantion/SB0/n3229 ), .C1(\U1/keyexpantion/SB0/n3246 ), .Y(
        \U1/keyexpantion/SB0/n1720 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1582  ( .A(
        \U1/keyexpantion/SB0/n3264 ), .B(\U1/keyexpantion/SB0/n3267 ), .Y(
        \U1/keyexpantion/SB0/n3050 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1581  ( .A(
        \U1/keyexpantion/SB0/n3252 ), .B(\U1/keyexpantion/SB0/n3194 ), .Y(
        \U1/keyexpantion/SB0/n3183 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1580  ( .A(
        \U1/keyexpantion/SB0/n3155 ), .B(\U1/keyexpantion/SB0/n3252 ), .Y(
        \U1/keyexpantion/SB0/n3117 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1579  ( .A(
        \U1/keyexpantion/SB0/n3139 ), .B(\U1/keyexpantion/SB0/n3219 ), .Y(
        \U1/keyexpantion/SB0/n2989 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1578  ( .AN(
        \U1/keyexpantion/SB0/n3050 ), .B(\U1/keyexpantion/SB0/n3183 ), .C(
        \U1/keyexpantion/SB0/n3117 ), .D(\U1/keyexpantion/SB0/n2989 ), .Y(
        \U1/keyexpantion/SB0/n1719 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1577  ( .A(
        \U1/keyexpantion/SB0/n3262 ), .B(\U1/keyexpantion/SB0/n3247 ), .Y(
        \U1/keyexpantion/SB0/n3062 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1576  ( .A(
        \U1/keyexpantion/SB0/n3139 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3129 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1575  ( .A(
        \U1/keyexpantion/SB0/n2991 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3030 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1574  ( .A(
        \U1/keyexpantion/SB0/n3198 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3075 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1573  ( .A(
        \U1/keyexpantion/SB0/n3062 ), .B(\U1/keyexpantion/SB0/n3129 ), .C(
        \U1/keyexpantion/SB0/n3030 ), .D(\U1/keyexpantion/SB0/n3075 ), .Y(
        \U1/keyexpantion/SB0/n1718 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1572  ( .A(\U1/keyexpantion/SB0/n1721 ), .B(\U1/keyexpantion/SB0/n1720 ), .C(\U1/keyexpantion/SB0/n1719 ), .D(
        \U1/keyexpantion/SB0/n1718 ), .Y(\U1/keyexpantion/SB0/n1722 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1571  ( .A(\U1/keyexpantion/SB0/n1722 ), .Y(\U1/keyexpantion/SB0/n3244 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1570  ( .A(
        \U1/keyexpantion/SB0/n3260 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n1723 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1569  ( .AN(
        \U1/keyexpantion/SB0/n2914 ), .B(\U1/keyexpantion/SB0/n1724 ), .C(
        \U1/keyexpantion/SB0/n3244 ), .D(\U1/keyexpantion/SB0/n1723 ), .Y(
        \U1/keyexpantion/SB0/n1725 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1568  ( .A(\U1/keyexpantion/SB0/n3023 ), .B(\U1/keyexpantion/SB0/n3120 ), .C(\U1/keyexpantion/SB0/n1728 ), .D(
        \U1/keyexpantion/SB0/n1727 ), .E(\U1/keyexpantion/SB0/n1726 ), .F(
        \U1/keyexpantion/SB0/n1725 ), .Y(\U1/keyexpantion/SB0/n2354 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1567  ( .A(
        \U1/keyexpantion/SB0/n3245 ), .B(\U1/keyexpantion/SB0/n2335 ), .Y(
        \U1/keyexpantion/SB0/n3068 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1566  ( .A(
        \U1/keyexpantion/SB0/n3195 ), .B(\U1/keyexpantion/SB0/n3262 ), .Y(
        \U1/keyexpantion/SB0/n3119 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1565  ( .A(
        \U1/keyexpantion/SB0/n3251 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3021 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1564  ( .A(\U1/keyexpantion/SB0/n2992 ), .Y(\U1/keyexpantion/SB0/n3240 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1563  ( .A(
        \U1/keyexpantion/SB0/n3240 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3044 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1562  ( .AN(
        \U1/keyexpantion/SB0/n3068 ), .B(\U1/keyexpantion/SB0/n3119 ), .C(
        \U1/keyexpantion/SB0/n3021 ), .D(\U1/keyexpantion/SB0/n3044 ), .Y(
        \U1/keyexpantion/SB0/n1735 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1561  ( .A(
        \U1/keyexpantion/SB0/n3232 ), .B(\U1/keyexpantion/SB0/n3103 ), .Y(
        \U1/keyexpantion/SB0/n3145 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1560  ( .A(
        \U1/keyexpantion/SB0/n3155 ), .B(\U1/keyexpantion/SB0/n3221 ), .Y(
        \U1/keyexpantion/SB0/n3001 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1559  ( .A0(
        \U1/keyexpantion/SB0/n3241 ), .A1(\U1/keyexpantion/SB0/n3161 ), .B0(
        \U1/keyexpantion/SB0/n2991 ), .Y(\U1/keyexpantion/SB0/n1729 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1558  ( .A(
        \U1/keyexpantion/SB0/n3222 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3093 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1557  ( .AN(
        \U1/keyexpantion/SB0/n3145 ), .B(\U1/keyexpantion/SB0/n3001 ), .C(
        \U1/keyexpantion/SB0/n1729 ), .D(\U1/keyexpantion/SB0/n3093 ), .Y(
        \U1/keyexpantion/SB0/n1730 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1556  ( .A(\U1/keyexpantion/SB0/n1730 ), .Y(\U1/keyexpantion/SB0/n1734 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1555  ( .A(\U1/keyexpantion/SB0/n3122 ), .Y(\U1/keyexpantion/SB0/n3242 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1554  ( .A(\U1/keyexpantion/SB0/n3267 ), .Y(\U1/keyexpantion/SB0/n3162 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1553  ( .A0(
        \U1/keyexpantion/SB0/n3262 ), .A1(\U1/keyexpantion/SB0/n3196 ), .B0(
        \U1/keyexpantion/SB0/n3242 ), .B1(\U1/keyexpantion/SB0/n3077 ), .C0(
        \U1/keyexpantion/SB0/n3162 ), .C1(\U1/keyexpantion/SB0/n3240 ), .Y(
        \U1/keyexpantion/SB0/n1733 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1552  ( .A0(
        \U1/keyexpantion/SB0/n3088 ), .A1(\U1/keyexpantion/SB0/n3245 ), .B0(
        \U1/keyexpantion/SB0/n3265 ), .B1(\U1/keyexpantion/SB0/n3266 ), .Y(
        \U1/keyexpantion/SB0/n1731 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1551  ( .A0(
        \U1/keyexpantion/SB0/n3139 ), .A1(\U1/keyexpantion/SB0/n2977 ), .B0(
        \U1/keyexpantion/SB0/n3195 ), .B1(\U1/keyexpantion/SB0/n3218 ), .C0(
        \U1/keyexpantion/SB0/n1731 ), .Y(\U1/keyexpantion/SB0/n1732 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1550  ( .AN(
        \U1/keyexpantion/SB0/n1735 ), .B(\U1/keyexpantion/SB0/n1734 ), .C(
        \U1/keyexpantion/SB0/n1733 ), .D(\U1/keyexpantion/SB0/n1732 ), .Y(
        \U1/keyexpantion/SB0/n2912 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1549  ( .A(
        \U1/keyexpantion/SB0/n3266 ), .B(\U1/keyexpantion/SB0/n3103 ), .Y(
        \U1/keyexpantion/SB0/n2986 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1548  ( .A0(
        \U1/keyexpantion/SB0/n3173 ), .A1(\U1/keyexpantion/SB0/n3266 ), .B0(
        \U1/keyexpantion/SB0/n3205 ), .Y(\U1/keyexpantion/SB0/n1740 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1547  ( .A(
        \U1/keyexpantion/SB0/n3205 ), .B(\U1/keyexpantion/SB0/n3193 ), .Y(
        \U1/keyexpantion/SB0/n3070 ) );
  AO22_X0P5M_A12TL \U1/keyexpantion/SB0/U1546  ( .A0(
        \U1/keyexpantion/SB0/n3194 ), .A1(\U1/keyexpantion/SB0/n2977 ), .B0(
        \U1/keyexpantion/SB0/n3070 ), .B1(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n1739 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1545  ( .A0(
        \U1/keyexpantion/SB0/n3227 ), .A1(\U1/keyexpantion/SB0/n3267 ), .B0(
        \U1/keyexpantion/SB0/n2992 ), .B1(\U1/keyexpantion/SB0/n3085 ), .C0(
        \U1/keyexpantion/SB0/n3229 ), .C1(\U1/keyexpantion/SB0/n3258 ), .Y(
        \U1/keyexpantion/SB0/n1738 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1544  ( .A(\U1/keyexpantion/SB0/n3088 ), .Y(\U1/keyexpantion/SB0/n3156 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1543  ( .A(
        \U1/keyexpantion/SB0/n3260 ), .B(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3182 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1542  ( .A(
        \U1/keyexpantion/SB0/n3155 ), .B(\U1/keyexpantion/SB0/n2977 ), .Y(
        \U1/keyexpantion/SB0/n3009 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1541  ( .A(
        \U1/keyexpantion/SB0/n2991 ), .B(\U1/keyexpantion/SB0/n3198 ), .Y(
        \U1/keyexpantion/SB0/n3029 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1540  ( .A(
        \U1/keyexpantion/SB0/n3155 ), .B(\U1/keyexpantion/SB0/n3196 ), .Y(
        \U1/keyexpantion/SB0/n3128 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1539  ( .A(
        \U1/keyexpantion/SB0/n3182 ), .B(\U1/keyexpantion/SB0/n3009 ), .C(
        \U1/keyexpantion/SB0/n3029 ), .D(\U1/keyexpantion/SB0/n3128 ), .Y(
        \U1/keyexpantion/SB0/n1737 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1538  ( .A(
        \U1/keyexpantion/SB0/n3175 ), .B(\U1/keyexpantion/SB0/n3088 ), .Y(
        \U1/keyexpantion/SB0/n3051 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1537  ( .A(
        \U1/keyexpantion/SB0/n3161 ), .B(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3061 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1536  ( .A(
        \U1/keyexpantion/SB0/n3222 ), .B(\U1/keyexpantion/SB0/n3077 ), .Y(
        \U1/keyexpantion/SB0/n3092 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1535  ( .AN(
        \U1/keyexpantion/SB0/n3051 ), .B(\U1/keyexpantion/SB0/n3061 ), .C(
        \U1/keyexpantion/SB0/n3092 ), .Y(\U1/keyexpantion/SB0/n1736 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1534  ( .A(\U1/keyexpantion/SB0/n2986 ), .B(\U1/keyexpantion/SB0/n1740 ), .C(\U1/keyexpantion/SB0/n1739 ), .D(
        \U1/keyexpantion/SB0/n1738 ), .E(\U1/keyexpantion/SB0/n1737 ), .F(
        \U1/keyexpantion/SB0/n1736 ), .Y(\U1/keyexpantion/SB0/n3273 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1533  ( .A0(
        \U1/keyexpantion/SB0/n2991 ), .A1(\U1/keyexpantion/SB0/n3219 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n1741 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1532  ( .A(
        \U1/keyexpantion/SB0/n2977 ), .B(\U1/keyexpantion/SB0/n3077 ), .Y(
        \U1/keyexpantion/SB0/n3114 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1531  ( .A(
        \U1/keyexpantion/SB0/n3194 ), .B(\U1/keyexpantion/SB0/n3242 ), .Y(
        \U1/keyexpantion/SB0/n3006 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1530  ( .A(
        \U1/keyexpantion/SB0/n3242 ), .B(\U1/keyexpantion/SB0/n3198 ), .Y(
        \U1/keyexpantion/SB0/n3057 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1529  ( .A(
        \U1/keyexpantion/SB0/n1741 ), .B(\U1/keyexpantion/SB0/n3114 ), .C(
        \U1/keyexpantion/SB0/n3006 ), .D(\U1/keyexpantion/SB0/n3057 ), .Y(
        \U1/keyexpantion/SB0/n1745 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1528  ( .A0(
        \U1/keyexpantion/SB0/n3245 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n2992 ), .B1(\U1/keyexpantion/SB0/n3217 ), .C0(
        \U1/keyexpantion/SB0/n3246 ), .C1(\U1/keyexpantion/SB0/n3103 ), .Y(
        \U1/keyexpantion/SB0/n1744 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1527  ( .A(
        \U1/keyexpantion/SB0/n3197 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3038 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1526  ( .A(
        \U1/keyexpantion/SB0/n3196 ), .B(\U1/keyexpantion/SB0/n3248 ), .Y(
        \U1/keyexpantion/SB0/n3178 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1525  ( .A(
        \U1/keyexpantion/SB0/n3196 ), .B(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3025 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1524  ( .A(
        \U1/keyexpantion/SB0/n3251 ), .B(\U1/keyexpantion/SB0/n3241 ), .Y(
        \U1/keyexpantion/SB0/n2987 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1523  ( .A(
        \U1/keyexpantion/SB0/n3038 ), .B(\U1/keyexpantion/SB0/n3178 ), .C(
        \U1/keyexpantion/SB0/n3025 ), .D(\U1/keyexpantion/SB0/n2987 ), .Y(
        \U1/keyexpantion/SB0/n1743 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1522  ( .A(
        \U1/keyexpantion/SB0/n3240 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3100 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1521  ( .A(
        \U1/keyexpantion/SB0/n3260 ), .B(\U1/keyexpantion/SB0/n3221 ), .Y(
        \U1/keyexpantion/SB0/n3073 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1520  ( .A(
        \U1/keyexpantion/SB0/n3250 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3124 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1519  ( .A(
        \U1/keyexpantion/SB0/n3003 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n2974 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1518  ( .A(
        \U1/keyexpantion/SB0/n3100 ), .B(\U1/keyexpantion/SB0/n3073 ), .C(
        \U1/keyexpantion/SB0/n3124 ), .D(\U1/keyexpantion/SB0/n2974 ), .Y(
        \U1/keyexpantion/SB0/n1742 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1517  ( .A(\U1/keyexpantion/SB0/n1745 ), .B(\U1/keyexpantion/SB0/n1744 ), .C(\U1/keyexpantion/SB0/n1743 ), .D(
        \U1/keyexpantion/SB0/n1742 ), .Y(\U1/keyexpantion/SB0/n2901 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1516  ( .A(\U1/keyexpantion/SB0/n2354 ), .B(\U1/keyexpantion/SB0/n2912 ), .C(\U1/keyexpantion/SB0/n3273 ), .D(
        \U1/keyexpantion/SB0/n2901 ), .Y(\U1/keyexpantion/SB0/n1755 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1515  ( .A(\U1/keyexpantion/SB0/n3227 ), .Y(\U1/keyexpantion/SB0/n3151 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1514  ( .A0(
        \U1/keyexpantion/SB0/n3103 ), .A1(\U1/keyexpantion/SB0/n2336 ), .B0(
        \U1/keyexpantion/SB0/n3072 ), .B1(\U1/keyexpantion/SB0/n3258 ), .Y(
        \U1/keyexpantion/SB0/n1746 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1513  ( .A0(
        \U1/keyexpantion/SB0/n3151 ), .A1(\U1/keyexpantion/SB0/n3203 ), .B0(
        \U1/keyexpantion/SB0/n3252 ), .B1(\U1/keyexpantion/SB0/n3260 ), .C0(
        \U1/keyexpantion/SB0/n1746 ), .Y(\U1/keyexpantion/SB0/n1754 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1512  ( .A(
        \U1/keyexpantion/SB0/n3172 ), .B(\U1/keyexpantion/SB0/n3175 ), .Y(
        \U1/keyexpantion/SB0/n3171 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1511  ( .A0(
        \U1/keyexpantion/SB0/n3106 ), .A1(\U1/keyexpantion/SB0/n3175 ), .B0(
        \U1/keyexpantion/SB0/n3088 ), .B1(\U1/keyexpantion/SB0/n3216 ), .Y(
        \U1/keyexpantion/SB0/n1747 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1510  ( .A0(
        \U1/keyexpantion/SB0/n3003 ), .A1(\U1/keyexpantion/SB0/n3171 ), .B0(
        \U1/keyexpantion/SB0/n3222 ), .B1(\U1/keyexpantion/SB0/n3241 ), .C0(
        \U1/keyexpantion/SB0/n1747 ), .Y(\U1/keyexpantion/SB0/n1753 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1509  ( .A(
        \U1/keyexpantion/SB0/n3246 ), .B(\U1/keyexpantion/SB0/n3105 ), .Y(
        \U1/keyexpantion/SB0/n1751 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1508  ( .A(
        \U1/keyexpantion/SB0/n3196 ), .B(\U1/keyexpantion/SB0/n3221 ), .Y(
        \U1/keyexpantion/SB0/n3163 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1507  ( .A(\U1/keyexpantion/SB0/n3163 ), .Y(\U1/keyexpantion/SB0/n1750 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1506  ( .A(
        \U1/keyexpantion/SB0/n3154 ), .B(\U1/keyexpantion/SB0/n3227 ), .Y(
        \U1/keyexpantion/SB0/n3035 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1505  ( .A(
        \U1/keyexpantion/SB0/n3232 ), .B(\U1/keyexpantion/SB0/n3230 ), .Y(
        \U1/keyexpantion/SB0/n3188 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1504  ( .A(\U1/keyexpantion/SB0/n3188 ), .Y(\U1/keyexpantion/SB0/n1748 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1503  ( .A(
        \U1/keyexpantion/SB0/n3203 ), .B(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3045 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1502  ( .AN(
        \U1/keyexpantion/SB0/n3035 ), .B(\U1/keyexpantion/SB0/n1748 ), .C(
        \U1/keyexpantion/SB0/n3045 ), .Y(\U1/keyexpantion/SB0/n1749 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1501  ( .A0(
        \U1/keyexpantion/SB0/n3162 ), .A1(\U1/keyexpantion/SB0/n1751 ), .B0(
        \U1/keyexpantion/SB0/n3139 ), .B1(\U1/keyexpantion/SB0/n1750 ), .C0(
        \U1/keyexpantion/SB0/n1749 ), .Y(\U1/keyexpantion/SB0/n1752 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1500  ( .AN(
        \U1/keyexpantion/SB0/n1755 ), .B(\U1/keyexpantion/SB0/n1754 ), .C(
        \U1/keyexpantion/SB0/n1753 ), .D(\U1/keyexpantion/SB0/n1752 ), .Y(
        \U1/keyexpantion/ws [0]) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1499  ( .A(\U1/rkey [6]), .Y(
        \U1/keyexpantion/SB0/n1762 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1498  ( .A(\U1/rkey [7]), .Y(
        \U1/keyexpantion/SB0/n1757 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1497  ( .A(
        \U1/keyexpantion/SB0/n1762 ), .B(\U1/keyexpantion/SB0/n1757 ), .Y(
        \U1/keyexpantion/SB0/n1767 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1496  ( .A(\U1/rkey [5]), .Y(
        \U1/keyexpantion/SB0/n1756 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1495  ( .A(
        \U1/keyexpantion/SB0/n1756 ), .B(\U1/rkey [4]), .Y(
        \U1/keyexpantion/SB0/n1774 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1494  ( .A(
        \U1/keyexpantion/SB0/n1767 ), .B(\U1/keyexpantion/SB0/n1774 ), .Y(
        \U1/keyexpantion/SB0/n3309 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1493  ( .A(\U1/rkey [3]), .Y(
        \U1/keyexpantion/SB0/n1765 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1492  ( .A(
        \U1/keyexpantion/SB0/n1765 ), .B(\U1/rkey [2]), .Y(
        \U1/keyexpantion/SB0/n1780 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1491  ( .A(\U1/rkey [0]), .Y(
        \U1/keyexpantion/SB0/n1758 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1490  ( .A(
        \U1/keyexpantion/SB0/n1758 ), .B(\U1/rkey [1]), .Y(
        \U1/keyexpantion/SB0/n1768 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1489  ( .A(
        \U1/keyexpantion/SB0/n1780 ), .B(\U1/keyexpantion/SB0/n1768 ), .Y(
        \U1/keyexpantion/SB0/n1919 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1488  ( .A(
        \U1/keyexpantion/SB0/n3309 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n1828 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1487  ( .A(\U1/rkey [1]), .Y(
        \U1/keyexpantion/SB0/n1759 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1486  ( .A(
        \U1/keyexpantion/SB0/n1759 ), .B(\U1/rkey [0]), .Y(
        \U1/keyexpantion/SB0/n1777 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1485  ( .A(\U1/rkey [2]), .Y(
        \U1/keyexpantion/SB0/n1764 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1484  ( .A(
        \U1/keyexpantion/SB0/n1764 ), .B(\U1/rkey [3]), .Y(
        \U1/keyexpantion/SB0/n1761 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1483  ( .A(
        \U1/keyexpantion/SB0/n1777 ), .B(\U1/keyexpantion/SB0/n1761 ), .Y(
        \U1/keyexpantion/SB0/n3355 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1482  ( .A(\U1/rkey [4]), .Y(
        \U1/keyexpantion/SB0/n1760 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1481  ( .A(
        \U1/keyexpantion/SB0/n1756 ), .B(\U1/keyexpantion/SB0/n1760 ), .Y(
        \U1/keyexpantion/SB0/n1788 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1480  ( .A(
        \U1/keyexpantion/SB0/n1757 ), .B(\U1/rkey [6]), .Y(
        \U1/keyexpantion/SB0/n1763 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1479  ( .A(
        \U1/keyexpantion/SB0/n1788 ), .B(\U1/keyexpantion/SB0/n1763 ), .Y(
        \U1/keyexpantion/SB0/n2028 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1478  ( .A0(
        \U1/keyexpantion/SB0/n1919 ), .A1(\U1/keyexpantion/SB0/n3355 ), .B0(
        \U1/keyexpantion/SB0/n2028 ), .Y(\U1/keyexpantion/SB0/n1773 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1477  ( .A(
        \U1/keyexpantion/SB0/n1759 ), .B(\U1/keyexpantion/SB0/n1758 ), .Y(
        \U1/keyexpantion/SB0/n1779 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1476  ( .A(
        \U1/keyexpantion/SB0/n1761 ), .B(\U1/keyexpantion/SB0/n1779 ), .Y(
        \U1/keyexpantion/SB0/n2027 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1475  ( .A(
        \U1/keyexpantion/SB0/n1760 ), .B(\U1/rkey [5]), .Y(
        \U1/keyexpantion/SB0/n1790 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1474  ( .A(
        \U1/keyexpantion/SB0/n1767 ), .B(\U1/keyexpantion/SB0/n1790 ), .Y(
        \U1/keyexpantion/SB0/n2002 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1473  ( .A(\U1/rkey [3]), .B(
        \U1/rkey [2]), .Y(\U1/keyexpantion/SB0/n1787 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1472  ( .A(
        \U1/keyexpantion/SB0/n1779 ), .B(\U1/keyexpantion/SB0/n1787 ), .Y(
        \U1/keyexpantion/SB0/n3310 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1471  ( .A(\U1/keyexpantion/SB0/n3310 ), .Y(\U1/keyexpantion/SB0/n3348 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1470  ( .A(\U1/rkey [1]), .B(
        \U1/rkey [0]), .Y(\U1/keyexpantion/SB0/n1786 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1469  ( .A(
        \U1/keyexpantion/SB0/n1761 ), .B(\U1/keyexpantion/SB0/n1786 ), .Y(
        \U1/keyexpantion/SB0/n3305 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1468  ( .A(\U1/keyexpantion/SB0/n3305 ), .Y(\U1/keyexpantion/SB0/n3342 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1467  ( .A(
        \U1/keyexpantion/SB0/n3348 ), .B(\U1/keyexpantion/SB0/n3342 ), .Y(
        \U1/keyexpantion/SB0/n1830 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1466  ( .A(\U1/rkey [7]), .B(
        \U1/rkey [6]), .Y(\U1/keyexpantion/SB0/n1781 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1465  ( .A(
        \U1/keyexpantion/SB0/n1774 ), .B(\U1/keyexpantion/SB0/n1781 ), .Y(
        \U1/keyexpantion/SB0/n3318 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1464  ( .A0(
        \U1/keyexpantion/SB0/n2027 ), .A1(\U1/keyexpantion/SB0/n2002 ), .B0(
        \U1/keyexpantion/SB0/n1830 ), .B1(\U1/keyexpantion/SB0/n3318 ), .Y(
        \U1/keyexpantion/SB0/n1772 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1463  ( .A(
        \U1/keyexpantion/SB0/n1761 ), .B(\U1/keyexpantion/SB0/n1768 ), .Y(
        \U1/keyexpantion/SB0/n1895 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1462  ( .A(
        \U1/keyexpantion/SB0/n1774 ), .B(\U1/keyexpantion/SB0/n1763 ), .Y(
        \U1/keyexpantion/SB0/n3353 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1461  ( .A(\U1/rkey [5]), .B(
        \U1/rkey [4]), .Y(\U1/keyexpantion/SB0/n1766 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1460  ( .A(
        \U1/keyexpantion/SB0/n1767 ), .B(\U1/keyexpantion/SB0/n1766 ), .Y(
        \U1/keyexpantion/SB0/n3289 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1459  ( .A(
        \U1/keyexpantion/SB0/n1790 ), .B(\U1/keyexpantion/SB0/n1763 ), .Y(
        \U1/keyexpantion/SB0/n3287 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1458  ( .A(
        \U1/keyexpantion/SB0/n1780 ), .B(\U1/keyexpantion/SB0/n1786 ), .Y(
        \U1/keyexpantion/SB0/n2017 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1457  ( .A0(
        \U1/keyexpantion/SB0/n1895 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n3310 ), .B1(\U1/keyexpantion/SB0/n3289 ), .C0(
        \U1/keyexpantion/SB0/n3287 ), .C1(\U1/keyexpantion/SB0/n2017 ), .Y(
        \U1/keyexpantion/SB0/n1771 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1456  ( .A(
        \U1/keyexpantion/SB0/n1762 ), .B(\U1/rkey [7]), .Y(
        \U1/keyexpantion/SB0/n1789 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1455  ( .A(
        \U1/keyexpantion/SB0/n1789 ), .B(\U1/keyexpantion/SB0/n1766 ), .Y(
        \U1/keyexpantion/SB0/n3317 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1454  ( .A(
        \U1/keyexpantion/SB0/n3317 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n1880 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1453  ( .A(
        \U1/keyexpantion/SB0/n1777 ), .B(\U1/keyexpantion/SB0/n1780 ), .Y(
        \U1/keyexpantion/SB0/n3351 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1452  ( .A(\U1/keyexpantion/SB0/n3351 ), .Y(\U1/keyexpantion/SB0/n2065 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1451  ( .A(
        \U1/keyexpantion/SB0/n1766 ), .B(\U1/keyexpantion/SB0/n1763 ), .Y(
        \U1/keyexpantion/SB0/n1813 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1450  ( .A(\U1/keyexpantion/SB0/n1813 ), .Y(\U1/keyexpantion/SB0/n3277 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1449  ( .A(
        \U1/keyexpantion/SB0/n2065 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n1863 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1448  ( .A(
        \U1/keyexpantion/SB0/n1765 ), .B(\U1/keyexpantion/SB0/n1764 ), .Y(
        \U1/keyexpantion/SB0/n1776 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1447  ( .A(
        \U1/keyexpantion/SB0/n1779 ), .B(\U1/keyexpantion/SB0/n1776 ), .Y(
        \U1/keyexpantion/SB0/n2013 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1446  ( .A(\U1/keyexpantion/SB0/n2013 ), .Y(\U1/keyexpantion/SB0/n2075 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U1445  ( .A(
        \U1/keyexpantion/SB0/n1781 ), .B(\U1/keyexpantion/SB0/n1766 ), .Y(
        \U1/keyexpantion/SB0/n3308 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1444  ( .A(
        \U1/keyexpantion/SB0/n2075 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1935 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1443  ( .A(
        \U1/keyexpantion/SB0/n1767 ), .B(\U1/keyexpantion/SB0/n1788 ), .Y(
        \U1/keyexpantion/SB0/n3356 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1442  ( .A(\U1/keyexpantion/SB0/n3356 ), .Y(\U1/keyexpantion/SB0/n3314 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1441  ( .A(
        \U1/keyexpantion/SB0/n3314 ), .B(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n1960 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1440  ( .AN(
        \U1/keyexpantion/SB0/n1880 ), .B(\U1/keyexpantion/SB0/n1863 ), .C(
        \U1/keyexpantion/SB0/n1935 ), .D(\U1/keyexpantion/SB0/n1960 ), .Y(
        \U1/keyexpantion/SB0/n1770 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1439  ( .A(\U1/keyexpantion/SB0/n2002 ), .Y(\U1/keyexpantion/SB0/n3278 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1438  ( .A(
        \U1/keyexpantion/SB0/n1787 ), .B(\U1/keyexpantion/SB0/n1768 ), .Y(
        \U1/keyexpantion/SB0/n2024 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1437  ( .A(\U1/keyexpantion/SB0/n2024 ), .Y(\U1/keyexpantion/SB0/n2061 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1436  ( .A(
        \U1/keyexpantion/SB0/n3278 ), .B(\U1/keyexpantion/SB0/n2061 ), .Y(
        \U1/keyexpantion/SB0/n1850 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1435  ( .A(\U1/keyexpantion/SB0/n3287 ), .Y(\U1/keyexpantion/SB0/n3341 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1434  ( .A(
        \U1/keyexpantion/SB0/n1768 ), .B(\U1/keyexpantion/SB0/n1776 ), .Y(
        \U1/keyexpantion/SB0/n2064 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1433  ( .A(\U1/keyexpantion/SB0/n2064 ), .Y(\U1/keyexpantion/SB0/n2026 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1432  ( .A(
        \U1/keyexpantion/SB0/n3341 ), .B(\U1/keyexpantion/SB0/n2026 ), .Y(
        \U1/keyexpantion/SB0/n1886 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1431  ( .A(
        \U1/keyexpantion/SB0/n3278 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1973 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U1430  ( .A(
        \U1/keyexpantion/SB0/n1850 ), .B(\U1/keyexpantion/SB0/n1886 ), .C(
        \U1/keyexpantion/SB0/n1973 ), .Y(\U1/keyexpantion/SB0/n1769 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1429  ( .A(\U1/keyexpantion/SB0/n1828 ), .B(\U1/keyexpantion/SB0/n1773 ), .C(\U1/keyexpantion/SB0/n1772 ), .D(
        \U1/keyexpantion/SB0/n1771 ), .E(\U1/keyexpantion/SB0/n1770 ), .F(
        \U1/keyexpantion/SB0/n1769 ), .Y(\U1/keyexpantion/SB0/n3362 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1428  ( .A(
        \U1/keyexpantion/SB0/n2002 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n1951 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1427  ( .A(\U1/keyexpantion/SB0/n2017 ), .Y(\U1/keyexpantion/SB0/n3339 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1426  ( .A(\U1/keyexpantion/SB0/n1895 ), .Y(\U1/keyexpantion/SB0/n3343 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1425  ( .A(
        \U1/keyexpantion/SB0/n1774 ), .B(\U1/keyexpantion/SB0/n1789 ), .Y(
        \U1/keyexpantion/SB0/n3352 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1424  ( .A(\U1/keyexpantion/SB0/n3352 ), .Y(\U1/keyexpantion/SB0/n3283 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1423  ( .A0(
        \U1/keyexpantion/SB0/n3339 ), .A1(\U1/keyexpantion/SB0/n3343 ), .B0(
        \U1/keyexpantion/SB0/n3283 ), .Y(\U1/keyexpantion/SB0/n1775 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1422  ( .A(
        \U1/keyexpantion/SB0/n3314 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1910 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1421  ( .A(\U1/keyexpantion/SB0/n2028 ), .Y(\U1/keyexpantion/SB0/n2060 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1420  ( .A(
        \U1/keyexpantion/SB0/n3348 ), .B(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n1872 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1419  ( .AN(
        \U1/keyexpantion/SB0/n1951 ), .B(\U1/keyexpantion/SB0/n1775 ), .C(
        \U1/keyexpantion/SB0/n1910 ), .D(\U1/keyexpantion/SB0/n1872 ), .Y(
        \U1/keyexpantion/SB0/n1785 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1418  ( .A(\U1/keyexpantion/SB0/n3318 ), .Y(\U1/keyexpantion/SB0/n1983 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1417  ( .A(
        \U1/keyexpantion/SB0/n1777 ), .B(\U1/keyexpantion/SB0/n1787 ), .Y(
        \U1/keyexpantion/SB0/n2046 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1416  ( .A(\U1/keyexpantion/SB0/n2046 ), .Y(\U1/keyexpantion/SB0/n3349 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1415  ( .A(\U1/keyexpantion/SB0/n3289 ), .Y(\U1/keyexpantion/SB0/n2062 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1414  ( .A(
        \U1/keyexpantion/SB0/n1786 ), .B(\U1/keyexpantion/SB0/n1776 ), .Y(
        \U1/keyexpantion/SB0/n3290 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1413  ( .A(\U1/keyexpantion/SB0/n3290 ), .Y(\U1/keyexpantion/SB0/n3340 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1412  ( .A0(
        \U1/keyexpantion/SB0/n1983 ), .A1(\U1/keyexpantion/SB0/n2075 ), .B0(
        \U1/keyexpantion/SB0/n3349 ), .B1(\U1/keyexpantion/SB0/n2062 ), .C0(
        \U1/keyexpantion/SB0/n3340 ), .C1(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n1784 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1411  ( .A(\U1/keyexpantion/SB0/n3309 ), .Y(\U1/keyexpantion/SB0/n1959 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1410  ( .A(
        \U1/keyexpantion/SB0/n1781 ), .B(\U1/keyexpantion/SB0/n1788 ), .Y(
        \U1/keyexpantion/SB0/n2077 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1409  ( .A(
        \U1/keyexpantion/SB0/n1777 ), .B(\U1/keyexpantion/SB0/n1776 ), .Y(
        \U1/keyexpantion/SB0/n3288 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1408  ( .A0(
        \U1/keyexpantion/SB0/n2077 ), .A1(\U1/keyexpantion/SB0/n3355 ), .B0(
        \U1/keyexpantion/SB0/n3288 ), .B1(\U1/keyexpantion/SB0/n2002 ), .Y(
        \U1/keyexpantion/SB0/n1778 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1407  ( .A0(
        \U1/keyexpantion/SB0/n2065 ), .A1(\U1/keyexpantion/SB0/n3314 ), .B0(
        \U1/keyexpantion/SB0/n1959 ), .B1(\U1/keyexpantion/SB0/n2026 ), .C0(
        \U1/keyexpantion/SB0/n1778 ), .Y(\U1/keyexpantion/SB0/n1783 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1406  ( .A(
        \U1/keyexpantion/SB0/n3277 ), .B(\U1/keyexpantion/SB0/n2026 ), .Y(
        \U1/keyexpantion/SB0/n1887 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1405  ( .A(
        \U1/keyexpantion/SB0/n1780 ), .B(\U1/keyexpantion/SB0/n1779 ), .Y(
        \U1/keyexpantion/SB0/n3311 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1404  ( .A(\U1/keyexpantion/SB0/n3311 ), .Y(\U1/keyexpantion/SB0/n3285 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1403  ( .A(
        \U1/keyexpantion/SB0/n3285 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n1852 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1402  ( .A(\U1/keyexpantion/SB0/n2077 ), .Y(\U1/keyexpantion/SB0/n3333 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1401  ( .A(
        \U1/keyexpantion/SB0/n3333 ), .B(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n1936 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1400  ( .A(
        \U1/keyexpantion/SB0/n1790 ), .B(\U1/keyexpantion/SB0/n1781 ), .Y(
        \U1/keyexpantion/SB0/n2072 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1399  ( .A(\U1/keyexpantion/SB0/n2072 ), .Y(\U1/keyexpantion/SB0/n3331 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1398  ( .A(
        \U1/keyexpantion/SB0/n3331 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1859 ) );
  AND4_X0P5M_A12TL \U1/keyexpantion/SB0/U1397  ( .A(
        \U1/keyexpantion/SB0/n1887 ), .B(\U1/keyexpantion/SB0/n1852 ), .C(
        \U1/keyexpantion/SB0/n1936 ), .D(\U1/keyexpantion/SB0/n1859 ), .Y(
        \U1/keyexpantion/SB0/n1782 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1396  ( .AN(
        \U1/keyexpantion/SB0/n1785 ), .B(\U1/keyexpantion/SB0/n1784 ), .C(
        \U1/keyexpantion/SB0/n1783 ), .D(\U1/keyexpantion/SB0/n1782 ), .Y(
        \U1/keyexpantion/SB0/n3304 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1395  ( .A(
        \U1/keyexpantion/SB0/n1787 ), .B(\U1/keyexpantion/SB0/n1786 ), .Y(
        \U1/keyexpantion/SB0/n3306 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1394  ( .A(
        \U1/keyexpantion/SB0/n3306 ), .B(\U1/keyexpantion/SB0/n2028 ), .Y(
        \U1/keyexpantion/SB0/n1972 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1393  ( .A(
        \U1/keyexpantion/SB0/n3309 ), .B(\U1/keyexpantion/SB0/n2013 ), .Y(
        \U1/keyexpantion/SB0/n1885 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1392  ( .A(
        \U1/keyexpantion/SB0/n3342 ), .B(\U1/keyexpantion/SB0/n3314 ), .Y(
        \U1/keyexpantion/SB0/n1849 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1391  ( .A0(
        \U1/keyexpantion/SB0/n3309 ), .A1(\U1/keyexpantion/SB0/n3351 ), .B0(
        \U1/keyexpantion/SB0/n1849 ), .Y(\U1/keyexpantion/SB0/n1794 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1390  ( .A(\U1/keyexpantion/SB0/n1919 ), .Y(\U1/keyexpantion/SB0/n3334 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1389  ( .A(
        \U1/keyexpantion/SB0/n3277 ), .B(\U1/keyexpantion/SB0/n3334 ), .Y(
        \U1/keyexpantion/SB0/n1984 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1388  ( .A(
        \U1/keyexpantion/SB0/n3277 ), .B(\U1/keyexpantion/SB0/n3343 ), .Y(
        \U1/keyexpantion/SB0/n1961 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1387  ( .A(
        \U1/keyexpantion/SB0/n1789 ), .B(\U1/keyexpantion/SB0/n1788 ), .Y(
        \U1/keyexpantion/SB0/n2015 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1386  ( .A(\U1/keyexpantion/SB0/n2015 ), .Y(\U1/keyexpantion/SB0/n3316 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1385  ( .A(
        \U1/keyexpantion/SB0/n3316 ), .B(\U1/keyexpantion/SB0/n2026 ), .Y(
        \U1/keyexpantion/SB0/n1862 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1384  ( .A(
        \U1/keyexpantion/SB0/n3316 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1909 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1383  ( .A(
        \U1/keyexpantion/SB0/n1984 ), .B(\U1/keyexpantion/SB0/n1961 ), .C(
        \U1/keyexpantion/SB0/n1862 ), .D(\U1/keyexpantion/SB0/n1909 ), .Y(
        \U1/keyexpantion/SB0/n1793 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1382  ( .A(\U1/keyexpantion/SB0/n3355 ), .Y(\U1/keyexpantion/SB0/n3284 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1381  ( .A(
        \U1/keyexpantion/SB0/n3284 ), .B(\U1/keyexpantion/SB0/n1983 ), .Y(
        \U1/keyexpantion/SB0/n1934 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1380  ( .A(\U1/keyexpantion/SB0/n3306 ), .Y(\U1/keyexpantion/SB0/n3291 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1379  ( .A(
        \U1/keyexpantion/SB0/n1983 ), .B(\U1/keyexpantion/SB0/n3291 ), .Y(
        \U1/keyexpantion/SB0/n1929 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1378  ( .A(
        \U1/keyexpantion/SB0/n3331 ), .B(\U1/keyexpantion/SB0/n3285 ), .Y(
        \U1/keyexpantion/SB0/n1837 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1377  ( .A(
        \U1/keyexpantion/SB0/n3308 ), .B(\U1/keyexpantion/SB0/n2026 ), .Y(
        \U1/keyexpantion/SB0/n1916 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1376  ( .A(
        \U1/keyexpantion/SB0/n1934 ), .B(\U1/keyexpantion/SB0/n1929 ), .C(
        \U1/keyexpantion/SB0/n1837 ), .D(\U1/keyexpantion/SB0/n1916 ), .Y(
        \U1/keyexpantion/SB0/n1792 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1375  ( .A(\U1/keyexpantion/SB0/n3288 ), .Y(\U1/keyexpantion/SB0/n3332 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1374  ( .A(
        \U1/keyexpantion/SB0/n3283 ), .B(\U1/keyexpantion/SB0/n3332 ), .Y(
        \U1/keyexpantion/SB0/n1827 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1373  ( .A(
        \U1/keyexpantion/SB0/n2061 ), .B(\U1/keyexpantion/SB0/n3283 ), .Y(
        \U1/keyexpantion/SB0/n1871 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1372  ( .A(
        \U1/keyexpantion/SB0/n1790 ), .B(\U1/keyexpantion/SB0/n1789 ), .Y(
        \U1/keyexpantion/SB0/n3312 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1371  ( .A(\U1/keyexpantion/SB0/n3312 ), .Y(\U1/keyexpantion/SB0/n3338 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1370  ( .A(
        \U1/keyexpantion/SB0/n2075 ), .B(\U1/keyexpantion/SB0/n3338 ), .Y(
        \U1/keyexpantion/SB0/n1897 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1369  ( .A(
        \U1/keyexpantion/SB0/n2061 ), .B(\U1/keyexpantion/SB0/n3333 ), .Y(
        \U1/keyexpantion/SB0/n1997 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1368  ( .A(
        \U1/keyexpantion/SB0/n1827 ), .B(\U1/keyexpantion/SB0/n1871 ), .C(
        \U1/keyexpantion/SB0/n1897 ), .D(\U1/keyexpantion/SB0/n1997 ), .Y(
        \U1/keyexpantion/SB0/n1791 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1367  ( .A(\U1/keyexpantion/SB0/n1972 ), .B(\U1/keyexpantion/SB0/n1885 ), .C(\U1/keyexpantion/SB0/n1794 ), .D(
        \U1/keyexpantion/SB0/n1793 ), .E(\U1/keyexpantion/SB0/n1792 ), .F(
        \U1/keyexpantion/SB0/n1791 ), .Y(\U1/keyexpantion/SB0/n3295 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1366  ( .A(
        \U1/keyexpantion/SB0/n3288 ), .B(\U1/keyexpantion/SB0/n2028 ), .Y(
        \U1/keyexpantion/SB0/n1838 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1365  ( .A(
        \U1/keyexpantion/SB0/n3289 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n1987 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1364  ( .A(
        \U1/keyexpantion/SB0/n3287 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n1879 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1363  ( .A(
        \U1/keyexpantion/SB0/n3287 ), .B(\U1/keyexpantion/SB0/n3290 ), .Y(
        \U1/keyexpantion/SB0/n1888 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1362  ( .A(
        \U1/keyexpantion/SB0/n3351 ), .B(\U1/keyexpantion/SB0/n3317 ), .Y(
        \U1/keyexpantion/SB0/n1926 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1361  ( .A(
        \U1/keyexpantion/SB0/n3316 ), .B(\U1/keyexpantion/SB0/n3334 ), .Y(
        \U1/keyexpantion/SB0/n1930 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1360  ( .A(
        \U1/keyexpantion/SB0/n2065 ), .B(\U1/keyexpantion/SB0/n3338 ), .Y(
        \U1/keyexpantion/SB0/n1851 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1359  ( .A(
        \U1/keyexpantion/SB0/n3340 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1864 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1358  ( .AN(
        \U1/keyexpantion/SB0/n1926 ), .B(\U1/keyexpantion/SB0/n1930 ), .C(
        \U1/keyexpantion/SB0/n1851 ), .D(\U1/keyexpantion/SB0/n1864 ), .Y(
        \U1/keyexpantion/SB0/n1798 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1357  ( .A(
        \U1/keyexpantion/SB0/n3309 ), .B(\U1/keyexpantion/SB0/n3290 ), .Y(
        \U1/keyexpantion/SB0/n1898 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1356  ( .A(
        \U1/keyexpantion/SB0/n3356 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n1974 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1355  ( .A(
        \U1/keyexpantion/SB0/n2002 ), .B(\U1/keyexpantion/SB0/n3355 ), .Y(
        \U1/keyexpantion/SB0/n1937 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1354  ( .A(
        \U1/keyexpantion/SB0/n2002 ), .B(\U1/keyexpantion/SB0/n2013 ), .Y(
        \U1/keyexpantion/SB0/n1835 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1353  ( .A0(
        \U1/keyexpantion/SB0/n3290 ), .A1(\U1/keyexpantion/SB0/n2002 ), .B0(
        \U1/keyexpantion/SB0/n3309 ), .B1(\U1/keyexpantion/SB0/n3355 ), .Y(
        \U1/keyexpantion/SB0/n1796 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1352  ( .A0(
        \U1/keyexpantion/SB0/n1895 ), .A1(\U1/keyexpantion/SB0/n2077 ), .B0(
        \U1/keyexpantion/SB0/n2027 ), .B1(\U1/keyexpantion/SB0/n3289 ), .Y(
        \U1/keyexpantion/SB0/n1795 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1351  ( .A(\U1/keyexpantion/SB0/n1898 ), .B(\U1/keyexpantion/SB0/n1974 ), .C(\U1/keyexpantion/SB0/n1937 ), .D(
        \U1/keyexpantion/SB0/n1835 ), .E(\U1/keyexpantion/SB0/n1796 ), .F(
        \U1/keyexpantion/SB0/n1795 ), .Y(\U1/keyexpantion/SB0/n1797 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1350  ( .A(\U1/keyexpantion/SB0/n1838 ), .B(\U1/keyexpantion/SB0/n1987 ), .C(\U1/keyexpantion/SB0/n1879 ), .D(
        \U1/keyexpantion/SB0/n1888 ), .E(\U1/keyexpantion/SB0/n1798 ), .F(
        \U1/keyexpantion/SB0/n1797 ), .Y(\U1/keyexpantion/SB0/n3330 ) );
  AOI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U1349  ( .A1N(
        \U1/keyexpantion/SB0/n3308 ), .A0(\U1/keyexpantion/SB0/n3352 ), .B0(
        \U1/keyexpantion/SB0/n2027 ), .Y(\U1/keyexpantion/SB0/n1799 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1348  ( .A(
        \U1/keyexpantion/SB0/n2002 ), .B(\U1/keyexpantion/SB0/n2046 ), .Y(
        \U1/keyexpantion/SB0/n1950 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1347  ( .A(
        \U1/keyexpantion/SB0/n3289 ), .B(\U1/keyexpantion/SB0/n2064 ), .Y(
        \U1/keyexpantion/SB0/n1857 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1346  ( .A(
        \U1/keyexpantion/SB0/n3289 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n1893 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1345  ( .A(\U1/keyexpantion/SB0/n1799 ), .B(\U1/keyexpantion/SB0/n1950 ), .C(\U1/keyexpantion/SB0/n1857 ), .D(
        \U1/keyexpantion/SB0/n1893 ), .Y(\U1/keyexpantion/SB0/n1804 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1344  ( .A0(
        \U1/keyexpantion/SB0/n2064 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n2028 ), .B1(\U1/keyexpantion/SB0/n3305 ), .C0(
        \U1/keyexpantion/SB0/n1919 ), .C1(\U1/keyexpantion/SB0/n3318 ), .Y(
        \U1/keyexpantion/SB0/n1803 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1343  ( .A(
        \U1/keyexpantion/SB0/n3351 ), .B(\U1/keyexpantion/SB0/n3318 ), .Y(
        \U1/keyexpantion/SB0/n1979 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1342  ( .A(
        \U1/keyexpantion/SB0/n2072 ), .B(\U1/keyexpantion/SB0/n2017 ), .Y(
        \U1/keyexpantion/SB0/n1840 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1341  ( .A(\U1/keyexpantion/SB0/n1840 ), .Y(\U1/keyexpantion/SB0/n1800 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1340  ( .A(
        \U1/keyexpantion/SB0/n3338 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1873 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1339  ( .A(
        \U1/keyexpantion/SB0/n1983 ), .B(\U1/keyexpantion/SB0/n2061 ), .Y(
        \U1/keyexpantion/SB0/n1860 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1338  ( .AN(
        \U1/keyexpantion/SB0/n1979 ), .B(\U1/keyexpantion/SB0/n1800 ), .C(
        \U1/keyexpantion/SB0/n1873 ), .D(\U1/keyexpantion/SB0/n1860 ), .Y(
        \U1/keyexpantion/SB0/n1802 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1337  ( .A(
        \U1/keyexpantion/SB0/n1895 ), .B(\U1/keyexpantion/SB0/n2028 ), .Y(
        \U1/keyexpantion/SB0/n1925 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1336  ( .A(
        \U1/keyexpantion/SB0/n1813 ), .B(\U1/keyexpantion/SB0/n3306 ), .Y(
        \U1/keyexpantion/SB0/n1902 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1335  ( .A(
        \U1/keyexpantion/SB0/n2015 ), .B(\U1/keyexpantion/SB0/n2027 ), .Y(
        \U1/keyexpantion/SB0/n1942 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1334  ( .A(
        \U1/keyexpantion/SB0/n2015 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n1834 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1333  ( .A(\U1/keyexpantion/SB0/n1925 ), .B(\U1/keyexpantion/SB0/n1902 ), .C(\U1/keyexpantion/SB0/n1942 ), .D(
        \U1/keyexpantion/SB0/n1834 ), .Y(\U1/keyexpantion/SB0/n1801 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1332  ( .A(\U1/keyexpantion/SB0/n1804 ), .B(\U1/keyexpantion/SB0/n1803 ), .C(\U1/keyexpantion/SB0/n1802 ), .D(
        \U1/keyexpantion/SB0/n1801 ), .Y(\U1/keyexpantion/SB0/n3302 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1331  ( .A(\U1/keyexpantion/SB0/n3317 ), .Y(\U1/keyexpantion/SB0/n3336 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1330  ( .A0(
        \U1/keyexpantion/SB0/n3339 ), .A1(\U1/keyexpantion/SB0/n3277 ), .B0(
        \U1/keyexpantion/SB0/n2075 ), .B1(\U1/keyexpantion/SB0/n3336 ), .Y(
        \U1/keyexpantion/SB0/n1805 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1329  ( .A0(
        \U1/keyexpantion/SB0/n3306 ), .A1(\U1/keyexpantion/SB0/n3356 ), .B0(
        \U1/keyexpantion/SB0/n3289 ), .B1(\U1/keyexpantion/SB0/n3355 ), .C0(
        \U1/keyexpantion/SB0/n1805 ), .Y(\U1/keyexpantion/SB0/n1811 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1328  ( .A(
        \U1/keyexpantion/SB0/n3312 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n1869 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1327  ( .A(
        \U1/keyexpantion/SB0/n3341 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1881 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1326  ( .A(
        \U1/keyexpantion/SB0/n3277 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1874 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1325  ( .A(
        \U1/keyexpantion/SB0/n3339 ), .B(\U1/keyexpantion/SB0/n3316 ), .Y(
        \U1/keyexpantion/SB0/n1846 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1324  ( .AN(
        \U1/keyexpantion/SB0/n1869 ), .B(\U1/keyexpantion/SB0/n1881 ), .C(
        \U1/keyexpantion/SB0/n1874 ), .D(\U1/keyexpantion/SB0/n1846 ), .Y(
        \U1/keyexpantion/SB0/n1810 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1323  ( .A(
        \U1/keyexpantion/SB0/n3290 ), .B(\U1/keyexpantion/SB0/n2064 ), .Y(
        \U1/keyexpantion/SB0/n1955 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1322  ( .A0(
        \U1/keyexpantion/SB0/n3334 ), .A1(\U1/keyexpantion/SB0/n1955 ), .B0(
        \U1/keyexpantion/SB0/n3331 ), .Y(\U1/keyexpantion/SB0/n1808 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1321  ( .A(\U1/keyexpantion/SB0/n3353 ), .Y(\U1/keyexpantion/SB0/n1956 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1320  ( .A0(
        \U1/keyexpantion/SB0/n2065 ), .A1(\U1/keyexpantion/SB0/n3332 ), .B0(
        \U1/keyexpantion/SB0/n1956 ), .Y(\U1/keyexpantion/SB0/n1807 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1319  ( .A(\U1/keyexpantion/SB0/n2027 ), .Y(\U1/keyexpantion/SB0/n2067 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1318  ( .A0(
        \U1/keyexpantion/SB0/n1959 ), .A1(\U1/keyexpantion/SB0/n1983 ), .B0(
        \U1/keyexpantion/SB0/n2067 ), .Y(\U1/keyexpantion/SB0/n1806 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1317  ( .A(
        \U1/keyexpantion/SB0/n2065 ), .B(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n1932 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1316  ( .A(
        \U1/keyexpantion/SB0/n1808 ), .B(\U1/keyexpantion/SB0/n1807 ), .C(
        \U1/keyexpantion/SB0/n1806 ), .D(\U1/keyexpantion/SB0/n1932 ), .Y(
        \U1/keyexpantion/SB0/n1809 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1315  ( .A(\U1/keyexpantion/SB0/n3295 ), .B(\U1/keyexpantion/SB0/n3330 ), .C(\U1/keyexpantion/SB0/n3302 ), .D(
        \U1/keyexpantion/SB0/n1811 ), .E(\U1/keyexpantion/SB0/n1810 ), .F(
        \U1/keyexpantion/SB0/n1809 ), .Y(\U1/keyexpantion/SB0/n2081 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1314  ( .A0(
        \U1/keyexpantion/SB0/n2026 ), .A1(\U1/keyexpantion/SB0/n3339 ), .B0(
        \U1/keyexpantion/SB0/n3333 ), .Y(\U1/keyexpantion/SB0/n1812 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1313  ( .A(
        \U1/keyexpantion/SB0/n3278 ), .B(\U1/keyexpantion/SB0/n2065 ), .Y(
        \U1/keyexpantion/SB0/n1917 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1312  ( .A(
        \U1/keyexpantion/SB0/n2062 ), .B(\U1/keyexpantion/SB0/n3285 ), .Y(
        \U1/keyexpantion/SB0/n1826 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1311  ( .A(
        \U1/keyexpantion/SB0/n3349 ), .B(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n1928 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1310  ( .A(
        \U1/keyexpantion/SB0/n1812 ), .B(\U1/keyexpantion/SB0/n1917 ), .C(
        \U1/keyexpantion/SB0/n1826 ), .D(\U1/keyexpantion/SB0/n1928 ), .Y(
        \U1/keyexpantion/SB0/n1817 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1309  ( .A0(
        \U1/keyexpantion/SB0/n2027 ), .A1(\U1/keyexpantion/SB0/n1813 ), .B0(
        \U1/keyexpantion/SB0/n3311 ), .B1(\U1/keyexpantion/SB0/n3356 ), .C0(
        \U1/keyexpantion/SB0/n3355 ), .C1(\U1/keyexpantion/SB0/n2072 ), .Y(
        \U1/keyexpantion/SB0/n1816 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1308  ( .A(
        \U1/keyexpantion/SB0/n1983 ), .B(\U1/keyexpantion/SB0/n3343 ), .Y(
        \U1/keyexpantion/SB0/n1848 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1307  ( .A(
        \U1/keyexpantion/SB0/n2065 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1971 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1306  ( .A(
        \U1/keyexpantion/SB0/n3284 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1870 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1305  ( .A(
        \U1/keyexpantion/SB0/n3349 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1933 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1304  ( .A(
        \U1/keyexpantion/SB0/n1848 ), .B(\U1/keyexpantion/SB0/n1971 ), .C(
        \U1/keyexpantion/SB0/n1870 ), .D(\U1/keyexpantion/SB0/n1933 ), .Y(
        \U1/keyexpantion/SB0/n1815 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1303  ( .A(
        \U1/keyexpantion/SB0/n3349 ), .B(\U1/keyexpantion/SB0/n3341 ), .Y(
        \U1/keyexpantion/SB0/n1896 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1302  ( .A(
        \U1/keyexpantion/SB0/n3342 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n1883 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1301  ( .A(
        \U1/keyexpantion/SB0/n3283 ), .B(\U1/keyexpantion/SB0/n3285 ), .Y(
        \U1/keyexpantion/SB0/n1861 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1300  ( .A(
        \U1/keyexpantion/SB0/n3332 ), .B(\U1/keyexpantion/SB0/n3336 ), .Y(
        \U1/keyexpantion/SB0/n1836 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1299  ( .A(
        \U1/keyexpantion/SB0/n1896 ), .B(\U1/keyexpantion/SB0/n1883 ), .C(
        \U1/keyexpantion/SB0/n1861 ), .D(\U1/keyexpantion/SB0/n1836 ), .Y(
        \U1/keyexpantion/SB0/n1814 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1298  ( .A(\U1/keyexpantion/SB0/n1817 ), .B(\U1/keyexpantion/SB0/n1816 ), .C(\U1/keyexpantion/SB0/n1815 ), .D(
        \U1/keyexpantion/SB0/n1814 ), .Y(\U1/keyexpantion/SB0/n1818 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1297  ( .A(\U1/keyexpantion/SB0/n1818 ), .Y(\U1/keyexpantion/SB0/n3293 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1296  ( .A0(
        \U1/keyexpantion/SB0/n3317 ), .A1(\U1/keyexpantion/SB0/n2046 ), .B0(
        \U1/keyexpantion/SB0/n3306 ), .B1(\U1/keyexpantion/SB0/n2077 ), .C0(
        \U1/keyexpantion/SB0/n3293 ), .Y(\U1/keyexpantion/SB0/n1825 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1295  ( .A(
        \U1/keyexpantion/SB0/n3338 ), .B(\U1/keyexpantion/SB0/n3283 ), .Y(
        \U1/keyexpantion/SB0/n1927 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U1294  ( .A1N(
        \U1/keyexpantion/SB0/n1927 ), .A0(\U1/keyexpantion/SB0/n3314 ), .B0(
        \U1/keyexpantion/SB0/n2026 ), .Y(\U1/keyexpantion/SB0/n1821 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1293  ( .A(
        \U1/keyexpantion/SB0/n2024 ), .B(\U1/keyexpantion/SB0/n3355 ), .Y(
        \U1/keyexpantion/SB0/n2025 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1292  ( .A0(
        \U1/keyexpantion/SB0/n3340 ), .A1(\U1/keyexpantion/SB0/n2025 ), .B0(
        \U1/keyexpantion/SB0/n3277 ), .Y(\U1/keyexpantion/SB0/n1820 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1291  ( .A0(
        \U1/keyexpantion/SB0/n2065 ), .A1(\U1/keyexpantion/SB0/n3342 ), .B0(
        \U1/keyexpantion/SB0/n2062 ), .Y(\U1/keyexpantion/SB0/n1819 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1290  ( .A(
        \U1/keyexpantion/SB0/n2061 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n1858 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1289  ( .A(
        \U1/keyexpantion/SB0/n1821 ), .B(\U1/keyexpantion/SB0/n1820 ), .C(
        \U1/keyexpantion/SB0/n1819 ), .D(\U1/keyexpantion/SB0/n1858 ), .Y(
        \U1/keyexpantion/SB0/n1824 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1288  ( .A(
        \U1/keyexpantion/SB0/n3284 ), .B(\U1/keyexpantion/SB0/n2067 ), .Y(
        \U1/keyexpantion/SB0/n2066 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1287  ( .A(
        \U1/keyexpantion/SB0/n2060 ), .B(\U1/keyexpantion/SB0/n1983 ), .Y(
        \U1/keyexpantion/SB0/n1822 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1286  ( .A0(
        \U1/keyexpantion/SB0/n2066 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n1822 ), .B1(\U1/keyexpantion/SB0/n2017 ), .C0(
        \U1/keyexpantion/SB0/n3311 ), .C1(\U1/keyexpantion/SB0/n3287 ), .Y(
        \U1/keyexpantion/SB0/n1823 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1285  ( .A(\U1/keyexpantion/SB0/n3362 ), .B(\U1/keyexpantion/SB0/n3304 ), .C(\U1/keyexpantion/SB0/n2081 ), .D(
        \U1/keyexpantion/SB0/n1825 ), .E(\U1/keyexpantion/SB0/n1824 ), .F(
        \U1/keyexpantion/SB0/n1823 ), .Y(\U1/keyexpantion/ws [10]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1284  ( .A(
        \U1/keyexpantion/SB0/n3356 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n2041 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1283  ( .A(
        \U1/keyexpantion/SB0/n3339 ), .B(\U1/keyexpantion/SB0/n1959 ), .Y(
        \U1/keyexpantion/SB0/n2043 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1282  ( .AN(
        \U1/keyexpantion/SB0/n1828 ), .B(\U1/keyexpantion/SB0/n1827 ), .C(
        \U1/keyexpantion/SB0/n1826 ), .D(\U1/keyexpantion/SB0/n2043 ), .Y(
        \U1/keyexpantion/SB0/n1833 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1281  ( .A(
        \U1/keyexpantion/SB0/n3333 ), .B(\U1/keyexpantion/SB0/n2062 ), .Y(
        \U1/keyexpantion/SB0/n1990 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1280  ( .A0(
        \U1/keyexpantion/SB0/n3278 ), .A1(\U1/keyexpantion/SB0/n3277 ), .B0(
        \U1/keyexpantion/SB0/n3332 ), .Y(\U1/keyexpantion/SB0/n1829 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1279  ( .A(
        \U1/keyexpantion/SB0/n3349 ), .B(\U1/keyexpantion/SB0/n1959 ), .Y(
        \U1/keyexpantion/SB0/n2068 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U1278  ( .A0(
        \U1/keyexpantion/SB0/n1990 ), .A1(\U1/keyexpantion/SB0/n3305 ), .B0(
        \U1/keyexpantion/SB0/n1829 ), .C0(\U1/keyexpantion/SB0/n2068 ), .Y(
        \U1/keyexpantion/SB0/n1832 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1277  ( .A0(
        \U1/keyexpantion/SB0/n2027 ), .A1(\U1/keyexpantion/SB0/n2077 ), .B0(
        \U1/keyexpantion/SB0/n1830 ), .B1(\U1/keyexpantion/SB0/n3317 ), .C0(
        \U1/keyexpantion/SB0/n3290 ), .C1(\U1/keyexpantion/SB0/n2072 ), .Y(
        \U1/keyexpantion/SB0/n1831 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1276  ( .A(\U1/keyexpantion/SB0/n1835 ), .B(\U1/keyexpantion/SB0/n2041 ), .C(\U1/keyexpantion/SB0/n1834 ), .D(
        \U1/keyexpantion/SB0/n1833 ), .E(\U1/keyexpantion/SB0/n1832 ), .F(
        \U1/keyexpantion/SB0/n1831 ), .Y(\U1/keyexpantion/SB0/n1969 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1275  ( .A(
        \U1/keyexpantion/SB0/n3332 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n2047 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1274  ( .AN(
        \U1/keyexpantion/SB0/n1838 ), .B(\U1/keyexpantion/SB0/n1837 ), .C(
        \U1/keyexpantion/SB0/n1836 ), .D(\U1/keyexpantion/SB0/n2047 ), .Y(
        \U1/keyexpantion/SB0/n1845 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1273  ( .A0(
        \U1/keyexpantion/SB0/n3340 ), .A1(\U1/keyexpantion/SB0/n3336 ), .B0(
        \U1/keyexpantion/SB0/n3341 ), .B1(\U1/keyexpantion/SB0/n3343 ), .C0(
        \U1/keyexpantion/SB0/n3283 ), .C1(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n1844 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1272  ( .A0(
        \U1/keyexpantion/SB0/n3310 ), .A1(\U1/keyexpantion/SB0/n3289 ), .B0(
        \U1/keyexpantion/SB0/n2028 ), .B1(\U1/keyexpantion/SB0/n2027 ), .Y(
        \U1/keyexpantion/SB0/n1839 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1271  ( .A0(
        \U1/keyexpantion/SB0/n1959 ), .A1(\U1/keyexpantion/SB0/n3332 ), .B0(
        \U1/keyexpantion/SB0/n3285 ), .B1(\U1/keyexpantion/SB0/n3308 ), .C0(
        \U1/keyexpantion/SB0/n1839 ), .Y(\U1/keyexpantion/SB0/n1843 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1270  ( .A(
        \U1/keyexpantion/SB0/n3317 ), .B(\U1/keyexpantion/SB0/n3352 ), .Y(
        \U1/keyexpantion/SB0/n3279 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1269  ( .A(
        \U1/keyexpantion/SB0/n3353 ), .B(\U1/keyexpantion/SB0/n3356 ), .Y(
        \U1/keyexpantion/SB0/n1841 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1268  ( .A0(
        \U1/keyexpantion/SB0/n3349 ), .A1(\U1/keyexpantion/SB0/n3279 ), .B0(
        \U1/keyexpantion/SB0/n2065 ), .B1(\U1/keyexpantion/SB0/n1841 ), .C0(
        \U1/keyexpantion/SB0/n1840 ), .Y(\U1/keyexpantion/SB0/n1842 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1267  ( .AN(
        \U1/keyexpantion/SB0/n1845 ), .B(\U1/keyexpantion/SB0/n1844 ), .C(
        \U1/keyexpantion/SB0/n1843 ), .D(\U1/keyexpantion/SB0/n1842 ), .Y(
        \U1/keyexpantion/SB0/n1995 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1266  ( .A(
        \U1/keyexpantion/SB0/n2002 ), .B(\U1/keyexpantion/SB0/n3311 ), .Y(
        \U1/keyexpantion/SB0/n2031 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1265  ( .A0(
        \U1/keyexpantion/SB0/n3312 ), .A1(\U1/keyexpantion/SB0/n3311 ), .B0(
        \U1/keyexpantion/SB0/n1846 ), .Y(\U1/keyexpantion/SB0/n1856 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1264  ( .A0(
        \U1/keyexpantion/SB0/n2065 ), .A1(\U1/keyexpantion/SB0/n3341 ), .B0(
        \U1/keyexpantion/SB0/n3284 ), .B1(\U1/keyexpantion/SB0/n3316 ), .Y(
        \U1/keyexpantion/SB0/n1847 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1263  ( .A0(
        \U1/keyexpantion/SB0/n3353 ), .A1(\U1/keyexpantion/SB0/n2046 ), .B0(
        \U1/keyexpantion/SB0/n2064 ), .B1(\U1/keyexpantion/SB0/n3352 ), .C0(
        \U1/keyexpantion/SB0/n1847 ), .Y(\U1/keyexpantion/SB0/n1855 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1262  ( .A(
        \U1/keyexpantion/SB0/n1919 ), .B(\U1/keyexpantion/SB0/n3317 ), .Y(
        \U1/keyexpantion/SB0/n3301 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1261  ( .A(
        \U1/keyexpantion/SB0/n3314 ), .B(\U1/keyexpantion/SB0/n3332 ), .Y(
        \U1/keyexpantion/SB0/n2044 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1260  ( .AN(
        \U1/keyexpantion/SB0/n3301 ), .B(\U1/keyexpantion/SB0/n1849 ), .C(
        \U1/keyexpantion/SB0/n1848 ), .D(\U1/keyexpantion/SB0/n2044 ), .Y(
        \U1/keyexpantion/SB0/n1854 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1259  ( .A(
        \U1/keyexpantion/SB0/n3289 ), .B(\U1/keyexpantion/SB0/n3306 ), .Y(
        \U1/keyexpantion/SB0/n2022 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1258  ( .AN(
        \U1/keyexpantion/SB0/n2022 ), .B(\U1/keyexpantion/SB0/n1852 ), .C(
        \U1/keyexpantion/SB0/n1851 ), .D(\U1/keyexpantion/SB0/n1850 ), .Y(
        \U1/keyexpantion/SB0/n1853 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1257  ( .A(\U1/keyexpantion/SB0/n2031 ), .B(\U1/keyexpantion/SB0/n1857 ), .C(\U1/keyexpantion/SB0/n1856 ), .D(
        \U1/keyexpantion/SB0/n1855 ), .E(\U1/keyexpantion/SB0/n1854 ), .F(
        \U1/keyexpantion/SB0/n1853 ), .Y(\U1/keyexpantion/SB0/n1931 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1256  ( .A(
        \U1/keyexpantion/SB0/n2024 ), .B(\U1/keyexpantion/SB0/n3309 ), .Y(
        \U1/keyexpantion/SB0/n2071 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1255  ( .A0(
        \U1/keyexpantion/SB0/n2024 ), .A1(\U1/keyexpantion/SB0/n3289 ), .B0(
        \U1/keyexpantion/SB0/n1858 ), .Y(\U1/keyexpantion/SB0/n1868 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1254  ( .A(
        \U1/keyexpantion/SB0/n3352 ), .B(\U1/keyexpantion/SB0/n1919 ), .Y(
        \U1/keyexpantion/SB0/n2030 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1253  ( .A(
        \U1/keyexpantion/SB0/n1956 ), .B(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n3321 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1252  ( .AN(
        \U1/keyexpantion/SB0/n2030 ), .B(\U1/keyexpantion/SB0/n1860 ), .C(
        \U1/keyexpantion/SB0/n1859 ), .D(\U1/keyexpantion/SB0/n3321 ), .Y(
        \U1/keyexpantion/SB0/n1867 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1251  ( .A(
        \U1/keyexpantion/SB0/n3283 ), .B(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n2052 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1250  ( .A(
        \U1/keyexpantion/SB0/n3348 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n3276 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1249  ( .A(
        \U1/keyexpantion/SB0/n2026 ), .B(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n3344 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1248  ( .A(
        \U1/keyexpantion/SB0/n1861 ), .B(\U1/keyexpantion/SB0/n2052 ), .C(
        \U1/keyexpantion/SB0/n3276 ), .D(\U1/keyexpantion/SB0/n3344 ), .Y(
        \U1/keyexpantion/SB0/n1866 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1247  ( .A(
        \U1/keyexpantion/SB0/n3331 ), .B(\U1/keyexpantion/SB0/n3342 ), .Y(
        \U1/keyexpantion/SB0/n2012 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1246  ( .A(
        \U1/keyexpantion/SB0/n1864 ), .B(\U1/keyexpantion/SB0/n1863 ), .C(
        \U1/keyexpantion/SB0/n2012 ), .D(\U1/keyexpantion/SB0/n1862 ), .Y(
        \U1/keyexpantion/SB0/n1865 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1245  ( .A(\U1/keyexpantion/SB0/n2071 ), .B(\U1/keyexpantion/SB0/n1869 ), .C(\U1/keyexpantion/SB0/n1868 ), .D(
        \U1/keyexpantion/SB0/n1867 ), .E(\U1/keyexpantion/SB0/n1866 ), .F(
        \U1/keyexpantion/SB0/n1865 ), .Y(\U1/keyexpantion/SB0/n1947 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1244  ( .A(
        \U1/keyexpantion/SB0/n3311 ), .B(\U1/keyexpantion/SB0/n2028 ), .Y(
        \U1/keyexpantion/SB0/n2023 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1243  ( .A(
        \U1/keyexpantion/SB0/n3333 ), .B(\U1/keyexpantion/SB0/n3340 ), .Y(
        \U1/keyexpantion/SB0/n2048 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1242  ( .A(
        \U1/keyexpantion/SB0/n3343 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n3274 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1241  ( .A(
        \U1/keyexpantion/SB0/n1871 ), .B(\U1/keyexpantion/SB0/n1870 ), .C(
        \U1/keyexpantion/SB0/n2048 ), .D(\U1/keyexpantion/SB0/n3274 ), .Y(
        \U1/keyexpantion/SB0/n1878 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1240  ( .A(
        \U1/keyexpantion/SB0/n1959 ), .B(\U1/keyexpantion/SB0/n3285 ), .Y(
        \U1/keyexpantion/SB0/n2034 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1239  ( .A(
        \U1/keyexpantion/SB0/n3342 ), .B(\U1/keyexpantion/SB0/n1959 ), .Y(
        \U1/keyexpantion/SB0/n3320 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1238  ( .A(
        \U1/keyexpantion/SB0/n1873 ), .B(\U1/keyexpantion/SB0/n2034 ), .C(
        \U1/keyexpantion/SB0/n1872 ), .D(\U1/keyexpantion/SB0/n3320 ), .Y(
        \U1/keyexpantion/SB0/n1877 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U1237  ( .A(
        \U1/keyexpantion/SB0/n2062 ), .B(\U1/keyexpantion/SB0/n3338 ), .C(
        \U1/keyexpantion/SB0/n2060 ), .Y(\U1/keyexpantion/SB0/n1875 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1236  ( .A0(
        \U1/keyexpantion/SB0/n1875 ), .A1(\U1/keyexpantion/SB0/n2017 ), .B0(
        \U1/keyexpantion/SB0/n2027 ), .B1(\U1/keyexpantion/SB0/n3356 ), .C0(
        \U1/keyexpantion/SB0/n1874 ), .Y(\U1/keyexpantion/SB0/n1876 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1235  ( .A(\U1/keyexpantion/SB0/n2023 ), .B(\U1/keyexpantion/SB0/n1880 ), .C(\U1/keyexpantion/SB0/n1879 ), .D(
        \U1/keyexpantion/SB0/n1878 ), .E(\U1/keyexpantion/SB0/n1877 ), .F(
        \U1/keyexpantion/SB0/n1876 ), .Y(\U1/keyexpantion/SB0/n1980 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1234  ( .A(
        \U1/keyexpantion/SB0/n3309 ), .B(\U1/keyexpantion/SB0/n1895 ), .Y(
        \U1/keyexpantion/SB0/n2035 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1233  ( .A0(
        \U1/keyexpantion/SB0/n2027 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n1881 ), .Y(\U1/keyexpantion/SB0/n1892 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1232  ( .A0(
        \U1/keyexpantion/SB0/n1983 ), .A1(\U1/keyexpantion/SB0/n2026 ), .B0(
        \U1/keyexpantion/SB0/n3331 ), .B1(\U1/keyexpantion/SB0/n3343 ), .Y(
        \U1/keyexpantion/SB0/n1882 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1231  ( .A0(
        \U1/keyexpantion/SB0/n3317 ), .A1(\U1/keyexpantion/SB0/n3355 ), .B0(
        \U1/keyexpantion/SB0/n3312 ), .B1(\U1/keyexpantion/SB0/n3288 ), .C0(
        \U1/keyexpantion/SB0/n1882 ), .Y(\U1/keyexpantion/SB0/n1891 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1230  ( .A(
        \U1/keyexpantion/SB0/n3312 ), .B(\U1/keyexpantion/SB0/n2027 ), .Y(
        \U1/keyexpantion/SB0/n3300 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1229  ( .A(\U1/keyexpantion/SB0/n3300 ), .Y(\U1/keyexpantion/SB0/n1884 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1228  ( .A(
        \U1/keyexpantion/SB0/n3341 ), .B(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n2054 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1227  ( .AN(
        \U1/keyexpantion/SB0/n1885 ), .B(\U1/keyexpantion/SB0/n1884 ), .C(
        \U1/keyexpantion/SB0/n1883 ), .D(\U1/keyexpantion/SB0/n2054 ), .Y(
        \U1/keyexpantion/SB0/n1890 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1226  ( .A(
        \U1/keyexpantion/SB0/n2065 ), .B(\U1/keyexpantion/SB0/n3316 ), .Y(
        \U1/keyexpantion/SB0/n2010 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1225  ( .AN(
        \U1/keyexpantion/SB0/n1888 ), .B(\U1/keyexpantion/SB0/n1887 ), .C(
        \U1/keyexpantion/SB0/n1886 ), .D(\U1/keyexpantion/SB0/n2010 ), .Y(
        \U1/keyexpantion/SB0/n1889 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1224  ( .A(\U1/keyexpantion/SB0/n2035 ), .B(\U1/keyexpantion/SB0/n1893 ), .C(\U1/keyexpantion/SB0/n1892 ), .D(
        \U1/keyexpantion/SB0/n1891 ), .E(\U1/keyexpantion/SB0/n1890 ), .F(
        \U1/keyexpantion/SB0/n1889 ), .Y(\U1/keyexpantion/SB0/n1954 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1223  ( .A0(
        \U1/keyexpantion/SB0/n2060 ), .A1(\U1/keyexpantion/SB0/n2025 ), .B0(
        \U1/keyexpantion/SB0/n1983 ), .B1(\U1/keyexpantion/SB0/n2067 ), .Y(
        \U1/keyexpantion/SB0/n1894 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1222  ( .A0(
        \U1/keyexpantion/SB0/n3290 ), .A1(\U1/keyexpantion/SB0/n3289 ), .B0(
        \U1/keyexpantion/SB0/n1895 ), .B1(\U1/keyexpantion/SB0/n3352 ), .C0(
        \U1/keyexpantion/SB0/n1894 ), .Y(\U1/keyexpantion/SB0/n1905 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1221  ( .A(
        \U1/keyexpantion/SB0/n3338 ), .B(\U1/keyexpantion/SB0/n3334 ), .Y(
        \U1/keyexpantion/SB0/n2051 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1220  ( .AN(
        \U1/keyexpantion/SB0/n1898 ), .B(\U1/keyexpantion/SB0/n1897 ), .C(
        \U1/keyexpantion/SB0/n1896 ), .D(\U1/keyexpantion/SB0/n2051 ), .Y(
        \U1/keyexpantion/SB0/n1904 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1219  ( .A0(
        \U1/keyexpantion/SB0/n3291 ), .A1(\U1/keyexpantion/SB0/n3349 ), .B0(
        \U1/keyexpantion/SB0/n3331 ), .Y(\U1/keyexpantion/SB0/n1901 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1218  ( .A(
        \U1/keyexpantion/SB0/n3353 ), .B(\U1/keyexpantion/SB0/n2002 ), .Y(
        \U1/keyexpantion/SB0/n1899 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1217  ( .A0(
        \U1/keyexpantion/SB0/n3342 ), .A1(\U1/keyexpantion/SB0/n1899 ), .B0(
        \U1/keyexpantion/SB0/n3338 ), .B1(\U1/keyexpantion/SB0/n1955 ), .Y(
        \U1/keyexpantion/SB0/n1900 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1216  ( .AN(
        \U1/keyexpantion/SB0/n1902 ), .B(\U1/keyexpantion/SB0/n1901 ), .C(
        \U1/keyexpantion/SB0/n1900 ), .Y(\U1/keyexpantion/SB0/n1903 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1215  ( .A(\U1/keyexpantion/SB0/n1947 ), .B(\U1/keyexpantion/SB0/n1980 ), .C(\U1/keyexpantion/SB0/n1954 ), .D(
        \U1/keyexpantion/SB0/n1905 ), .E(\U1/keyexpantion/SB0/n1904 ), .F(
        \U1/keyexpantion/SB0/n1903 ), .Y(\U1/keyexpantion/SB0/n2006 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1214  ( .A(\U1/keyexpantion/SB0/n1969 ), .B(\U1/keyexpantion/SB0/n1995 ), .C(\U1/keyexpantion/SB0/n1931 ), .D(
        \U1/keyexpantion/SB0/n2006 ), .Y(\U1/keyexpantion/SB0/n1915 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1213  ( .A(
        \U1/keyexpantion/SB0/n3342 ), .B(\U1/keyexpantion/SB0/n2075 ), .Y(
        \U1/keyexpantion/SB0/n2016 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1212  ( .A(
        \U1/keyexpantion/SB0/n3332 ), .B(\U1/keyexpantion/SB0/n2067 ), .Y(
        \U1/keyexpantion/SB0/n2009 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1211  ( .A(
        \U1/keyexpantion/SB0/n3306 ), .B(\U1/keyexpantion/SB0/n3311 ), .Y(
        \U1/keyexpantion/SB0/n3315 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1210  ( .A0(
        \U1/keyexpantion/SB0/n1959 ), .A1(\U1/keyexpantion/SB0/n3284 ), .B0(
        \U1/keyexpantion/SB0/n3315 ), .B1(\U1/keyexpantion/SB0/n3314 ), .Y(
        \U1/keyexpantion/SB0/n1906 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1209  ( .A0(
        \U1/keyexpantion/SB0/n2028 ), .A1(\U1/keyexpantion/SB0/n2016 ), .B0(
        \U1/keyexpantion/SB0/n3287 ), .B1(\U1/keyexpantion/SB0/n2009 ), .C0(
        \U1/keyexpantion/SB0/n1906 ), .Y(\U1/keyexpantion/SB0/n1907 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1208  ( .A(\U1/keyexpantion/SB0/n1907 ), .Y(\U1/keyexpantion/SB0/n1914 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1207  ( .A0(
        \U1/keyexpantion/SB0/n3310 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n2027 ), .B1(\U1/keyexpantion/SB0/n2002 ), .Y(
        \U1/keyexpantion/SB0/n1908 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1206  ( .A0(
        \U1/keyexpantion/SB0/n2061 ), .A1(\U1/keyexpantion/SB0/n3277 ), .B0(
        \U1/keyexpantion/SB0/n3336 ), .B1(\U1/keyexpantion/SB0/n3291 ), .C0(
        \U1/keyexpantion/SB0/n1908 ), .Y(\U1/keyexpantion/SB0/n1913 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1205  ( .A0(
        \U1/keyexpantion/SB0/n2075 ), .A1(\U1/keyexpantion/SB0/n3332 ), .B0(
        \U1/keyexpantion/SB0/n2062 ), .Y(\U1/keyexpantion/SB0/n1911 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1204  ( .A(
        \U1/keyexpantion/SB0/n3349 ), .B(\U1/keyexpantion/SB0/n3314 ), .Y(
        \U1/keyexpantion/SB0/n2033 ) );
  AND4_X0P5M_A12TL \U1/keyexpantion/SB0/U1203  ( .A(
        \U1/keyexpantion/SB0/n1911 ), .B(\U1/keyexpantion/SB0/n2033 ), .C(
        \U1/keyexpantion/SB0/n1910 ), .D(\U1/keyexpantion/SB0/n1909 ), .Y(
        \U1/keyexpantion/SB0/n1912 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1202  ( .AN(
        \U1/keyexpantion/SB0/n1915 ), .B(\U1/keyexpantion/SB0/n1914 ), .C(
        \U1/keyexpantion/SB0/n1913 ), .D(\U1/keyexpantion/SB0/n1912 ), .Y(
        \U1/keyexpantion/ws [11]) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1201  ( .A0(
        \U1/keyexpantion/SB0/n1927 ), .A1(\U1/keyexpantion/SB0/n2015 ), .B0(
        \U1/keyexpantion/SB0/n3306 ), .Y(\U1/keyexpantion/SB0/n1924 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1200  ( .A(
        \U1/keyexpantion/SB0/n1956 ), .B(\U1/keyexpantion/SB0/n3334 ), .Y(
        \U1/keyexpantion/SB0/n2042 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U1199  ( .A(
        \U1/keyexpantion/SB0/n1917 ), .B(\U1/keyexpantion/SB0/n2042 ), .C(
        \U1/keyexpantion/SB0/n1916 ), .Y(\U1/keyexpantion/SB0/n1923 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1198  ( .A(
        \U1/keyexpantion/SB0/n2060 ), .B(\U1/keyexpantion/SB0/n3331 ), .Y(
        \U1/keyexpantion/SB0/n1920 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1197  ( .A(
        \U1/keyexpantion/SB0/n3314 ), .B(\U1/keyexpantion/SB0/n1959 ), .Y(
        \U1/keyexpantion/SB0/n1918 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1196  ( .A0(
        \U1/keyexpantion/SB0/n1920 ), .A1(\U1/keyexpantion/SB0/n1919 ), .B0(
        \U1/keyexpantion/SB0/n1918 ), .B1(\U1/keyexpantion/SB0/n2064 ), .C0(
        \U1/keyexpantion/SB0/n2013 ), .C1(\U1/keyexpantion/SB0/n2015 ), .Y(
        \U1/keyexpantion/SB0/n1922 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1195  ( .A0(
        \U1/keyexpantion/SB0/n3312 ), .A1(\U1/keyexpantion/SB0/n2024 ), .B0(
        \U1/keyexpantion/SB0/n3290 ), .B1(\U1/keyexpantion/SB0/n3352 ), .C0(
        \U1/keyexpantion/SB0/n3317 ), .C1(\U1/keyexpantion/SB0/n2017 ), .Y(
        \U1/keyexpantion/SB0/n1921 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1194  ( .A(\U1/keyexpantion/SB0/n1926 ), .B(\U1/keyexpantion/SB0/n1925 ), .C(\U1/keyexpantion/SB0/n1924 ), .D(
        \U1/keyexpantion/SB0/n1923 ), .E(\U1/keyexpantion/SB0/n1922 ), .F(
        \U1/keyexpantion/SB0/n1921 ), .Y(\U1/keyexpantion/SB0/n2007 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1193  ( .A0(
        \U1/keyexpantion/SB0/n1927 ), .A1(\U1/keyexpantion/SB0/n3289 ), .B0(
        \U1/keyexpantion/SB0/n3355 ), .Y(\U1/keyexpantion/SB0/n1953 ) );
  AOI31_X0P5M_A12TL \U1/keyexpantion/SB0/U1192  ( .A0(
        \U1/keyexpantion/SB0/n3305 ), .A1(\U1/keyexpantion/SB0/n3288 ), .A2(
        \U1/keyexpantion/SB0/n2017 ), .B0(\U1/keyexpantion/SB0/n3318 ), .Y(
        \U1/keyexpantion/SB0/n1952 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1191  ( .A(
        \U1/keyexpantion/SB0/n3285 ), .B(\U1/keyexpantion/SB0/n3336 ), .Y(
        \U1/keyexpantion/SB0/n2049 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1190  ( .A(
        \U1/keyexpantion/SB0/n1930 ), .B(\U1/keyexpantion/SB0/n1929 ), .C(
        \U1/keyexpantion/SB0/n1928 ), .D(\U1/keyexpantion/SB0/n2049 ), .Y(
        \U1/keyexpantion/SB0/n1949 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1189  ( .A(\U1/keyexpantion/SB0/n1931 ), .Y(\U1/keyexpantion/SB0/n1946 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1188  ( .A(
        \U1/keyexpantion/SB0/n3318 ), .B(\U1/keyexpantion/SB0/n3311 ), .Y(
        \U1/keyexpantion/SB0/n2029 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1187  ( .A0(
        \U1/keyexpantion/SB0/n2009 ), .A1(\U1/keyexpantion/SB0/n2072 ), .B0(
        \U1/keyexpantion/SB0/n1932 ), .Y(\U1/keyexpantion/SB0/n1941 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1186  ( .A0(
        \U1/keyexpantion/SB0/n3289 ), .A1(\U1/keyexpantion/SB0/n3351 ), .B0(
        \U1/keyexpantion/SB0/n3306 ), .B1(\U1/keyexpantion/SB0/n2002 ), .C0(
        \U1/keyexpantion/SB0/n3290 ), .C1(\U1/keyexpantion/SB0/n3318 ), .Y(
        \U1/keyexpantion/SB0/n1940 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1185  ( .A(
        \U1/keyexpantion/SB0/n3316 ), .B(\U1/keyexpantion/SB0/n3332 ), .Y(
        \U1/keyexpantion/SB0/n2053 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1184  ( .A(
        \U1/keyexpantion/SB0/n2075 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n3281 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1183  ( .A(
        \U1/keyexpantion/SB0/n1934 ), .B(\U1/keyexpantion/SB0/n1933 ), .C(
        \U1/keyexpantion/SB0/n2053 ), .D(\U1/keyexpantion/SB0/n3281 ), .Y(
        \U1/keyexpantion/SB0/n1939 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1182  ( .A(
        \U1/keyexpantion/SB0/n3342 ), .B(\U1/keyexpantion/SB0/n3308 ), .Y(
        \U1/keyexpantion/SB0/n2011 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1181  ( .AN(
        \U1/keyexpantion/SB0/n1937 ), .B(\U1/keyexpantion/SB0/n1936 ), .C(
        \U1/keyexpantion/SB0/n1935 ), .D(\U1/keyexpantion/SB0/n2011 ), .Y(
        \U1/keyexpantion/SB0/n1938 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1180  ( .A(\U1/keyexpantion/SB0/n2029 ), .B(\U1/keyexpantion/SB0/n1942 ), .C(\U1/keyexpantion/SB0/n1941 ), .D(
        \U1/keyexpantion/SB0/n1940 ), .E(\U1/keyexpantion/SB0/n1939 ), .F(
        \U1/keyexpantion/SB0/n1938 ), .Y(\U1/keyexpantion/SB0/n1943 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1179  ( .A(\U1/keyexpantion/SB0/n1943 ), .Y(\U1/keyexpantion/SB0/n1996 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1178  ( .A0(
        \U1/keyexpantion/SB0/n3353 ), .A1(\U1/keyexpantion/SB0/n2024 ), .B0(
        \U1/keyexpantion/SB0/n3290 ), .B1(\U1/keyexpantion/SB0/n3356 ), .Y(
        \U1/keyexpantion/SB0/n1944 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1177  ( .A0(
        \U1/keyexpantion/SB0/n3333 ), .A1(\U1/keyexpantion/SB0/n3332 ), .B0(
        \U1/keyexpantion/SB0/n3339 ), .B1(\U1/keyexpantion/SB0/n3308 ), .C0(
        \U1/keyexpantion/SB0/n1944 ), .Y(\U1/keyexpantion/SB0/n1945 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1176  ( .AN(
        \U1/keyexpantion/SB0/n1947 ), .B(\U1/keyexpantion/SB0/n1946 ), .C(
        \U1/keyexpantion/SB0/n1996 ), .D(\U1/keyexpantion/SB0/n1945 ), .Y(
        \U1/keyexpantion/SB0/n1948 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1175  ( .A(\U1/keyexpantion/SB0/n1953 ), .B(\U1/keyexpantion/SB0/n1952 ), .C(\U1/keyexpantion/SB0/n1951 ), .D(
        \U1/keyexpantion/SB0/n1950 ), .E(\U1/keyexpantion/SB0/n1949 ), .F(
        \U1/keyexpantion/SB0/n1948 ), .Y(\U1/keyexpantion/SB0/n1994 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1174  ( .A(\U1/keyexpantion/SB0/n1954 ), .Y(\U1/keyexpantion/SB0/n1958 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1173  ( .A0(
        \U1/keyexpantion/SB0/n1956 ), .A1(\U1/keyexpantion/SB0/n1955 ), .B0(
        \U1/keyexpantion/SB0/n1959 ), .B1(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n1957 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U1172  ( .A0(
        \U1/keyexpantion/SB0/n2013 ), .A1(\U1/keyexpantion/SB0/n3318 ), .B0(
        \U1/keyexpantion/SB0/n1958 ), .C0(\U1/keyexpantion/SB0/n1957 ), .Y(
        \U1/keyexpantion/SB0/n1968 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1171  ( .A0(
        \U1/keyexpantion/SB0/n3285 ), .A1(\U1/keyexpantion/SB0/n3284 ), .B0(
        \U1/keyexpantion/SB0/n3341 ), .Y(\U1/keyexpantion/SB0/n1963 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1170  ( .A0(
        \U1/keyexpantion/SB0/n1959 ), .A1(\U1/keyexpantion/SB0/n3277 ), .B0(
        \U1/keyexpantion/SB0/n2067 ), .Y(\U1/keyexpantion/SB0/n1962 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1169  ( .A(
        \U1/keyexpantion/SB0/n1963 ), .B(\U1/keyexpantion/SB0/n1962 ), .C(
        \U1/keyexpantion/SB0/n1961 ), .D(\U1/keyexpantion/SB0/n1960 ), .Y(
        \U1/keyexpantion/SB0/n1967 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1168  ( .A(
        \U1/keyexpantion/SB0/n3334 ), .B(\U1/keyexpantion/SB0/n3343 ), .Y(
        \U1/keyexpantion/SB0/n1965 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1167  ( .A(
        \U1/keyexpantion/SB0/n3340 ), .B(\U1/keyexpantion/SB0/n3342 ), .Y(
        \U1/keyexpantion/SB0/n1964 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1166  ( .A(
        \U1/keyexpantion/SB0/n1983 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n3319 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1165  ( .A0(
        \U1/keyexpantion/SB0/n1965 ), .A1(\U1/keyexpantion/SB0/n2077 ), .B0(
        \U1/keyexpantion/SB0/n1964 ), .B1(\U1/keyexpantion/SB0/n2015 ), .C0(
        \U1/keyexpantion/SB0/n3319 ), .C1(\U1/keyexpantion/SB0/n2046 ), .Y(
        \U1/keyexpantion/SB0/n1966 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1164  ( .A(\U1/keyexpantion/SB0/n2007 ), .B(\U1/keyexpantion/SB0/n1994 ), .C(\U1/keyexpantion/SB0/n1969 ), .D(
        \U1/keyexpantion/SB0/n1968 ), .E(\U1/keyexpantion/SB0/n1967 ), .F(
        \U1/keyexpantion/SB0/n1966 ), .Y(\U1/keyexpantion/ws [12]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1163  ( .A(
        \U1/keyexpantion/SB0/n3309 ), .B(\U1/keyexpantion/SB0/n3306 ), .Y(
        \U1/keyexpantion/SB0/n2032 ) );
  AOI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U1162  ( .A1N(
        \U1/keyexpantion/SB0/n3315 ), .A0(\U1/keyexpantion/SB0/n3288 ), .B0(
        \U1/keyexpantion/SB0/n3353 ), .Y(\U1/keyexpantion/SB0/n1978 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1161  ( .A(
        \U1/keyexpantion/SB0/n2060 ), .B(\U1/keyexpantion/SB0/n3277 ), .Y(
        \U1/keyexpantion/SB0/n1970 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1160  ( .A0(
        \U1/keyexpantion/SB0/n2077 ), .A1(\U1/keyexpantion/SB0/n3311 ), .B0(
        \U1/keyexpantion/SB0/n1970 ), .B1(\U1/keyexpantion/SB0/n3290 ), .C0(
        \U1/keyexpantion/SB0/n3306 ), .C1(\U1/keyexpantion/SB0/n3287 ), .Y(
        \U1/keyexpantion/SB0/n1977 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1159  ( .A(
        \U1/keyexpantion/SB0/n3336 ), .B(\U1/keyexpantion/SB0/n2026 ), .Y(
        \U1/keyexpantion/SB0/n2050 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1158  ( .A(
        \U1/keyexpantion/SB0/n3308 ), .B(\U1/keyexpantion/SB0/n3291 ), .Y(
        \U1/keyexpantion/SB0/n3275 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1157  ( .AN(
        \U1/keyexpantion/SB0/n1972 ), .B(\U1/keyexpantion/SB0/n1971 ), .C(
        \U1/keyexpantion/SB0/n2050 ), .D(\U1/keyexpantion/SB0/n3275 ), .Y(
        \U1/keyexpantion/SB0/n1976 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1156  ( .A(
        \U1/keyexpantion/SB0/n3278 ), .B(\U1/keyexpantion/SB0/n3339 ), .Y(
        \U1/keyexpantion/SB0/n3322 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1155  ( .AN(
        \U1/keyexpantion/SB0/n1974 ), .B(\U1/keyexpantion/SB0/n1973 ), .C(
        \U1/keyexpantion/SB0/n3322 ), .Y(\U1/keyexpantion/SB0/n1975 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1154  ( .A(\U1/keyexpantion/SB0/n2032 ), .B(\U1/keyexpantion/SB0/n1979 ), .C(\U1/keyexpantion/SB0/n1978 ), .D(
        \U1/keyexpantion/SB0/n1977 ), .E(\U1/keyexpantion/SB0/n1976 ), .F(
        \U1/keyexpantion/SB0/n1975 ), .Y(\U1/keyexpantion/SB0/n2008 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1153  ( .A(\U1/keyexpantion/SB0/n1980 ), .Y(\U1/keyexpantion/SB0/n1982 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1152  ( .A0(
        \U1/keyexpantion/SB0/n3331 ), .A1(\U1/keyexpantion/SB0/n2065 ), .B0(
        \U1/keyexpantion/SB0/n2067 ), .B1(\U1/keyexpantion/SB0/n3336 ), .Y(
        \U1/keyexpantion/SB0/n1981 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U1151  ( .A0(
        \U1/keyexpantion/SB0/n3353 ), .A1(\U1/keyexpantion/SB0/n3355 ), .B0(
        \U1/keyexpantion/SB0/n1982 ), .C0(\U1/keyexpantion/SB0/n1981 ), .Y(
        \U1/keyexpantion/SB0/n1993 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1150  ( .A0(
        \U1/keyexpantion/SB0/n3333 ), .A1(\U1/keyexpantion/SB0/n3331 ), .B0(
        \U1/keyexpantion/SB0/n2026 ), .Y(\U1/keyexpantion/SB0/n1986 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1149  ( .A0(
        \U1/keyexpantion/SB0/n3334 ), .A1(\U1/keyexpantion/SB0/n3348 ), .B0(
        \U1/keyexpantion/SB0/n1983 ), .Y(\U1/keyexpantion/SB0/n1985 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1148  ( .AN(
        \U1/keyexpantion/SB0/n1987 ), .B(\U1/keyexpantion/SB0/n1986 ), .C(
        \U1/keyexpantion/SB0/n1985 ), .D(\U1/keyexpantion/SB0/n1984 ), .Y(
        \U1/keyexpantion/SB0/n1992 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1147  ( .A0(
        \U1/keyexpantion/SB0/n3341 ), .A1(\U1/keyexpantion/SB0/n3338 ), .B0(
        \U1/keyexpantion/SB0/n3342 ), .Y(\U1/keyexpantion/SB0/n1989 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1146  ( .A(
        \U1/keyexpantion/SB0/n2024 ), .B(\U1/keyexpantion/SB0/n3311 ), .Y(
        \U1/keyexpantion/SB0/n3350 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1145  ( .A0(
        \U1/keyexpantion/SB0/n3316 ), .A1(\U1/keyexpantion/SB0/n3350 ), .B0(
        \U1/keyexpantion/SB0/n2061 ), .B1(\U1/keyexpantion/SB0/n3314 ), .Y(
        \U1/keyexpantion/SB0/n1988 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U1144  ( .A0(
        \U1/keyexpantion/SB0/n1990 ), .A1(\U1/keyexpantion/SB0/n2046 ), .B0(
        \U1/keyexpantion/SB0/n1989 ), .C0(\U1/keyexpantion/SB0/n1988 ), .Y(
        \U1/keyexpantion/SB0/n1991 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1143  ( .A(\U1/keyexpantion/SB0/n2008 ), .B(\U1/keyexpantion/SB0/n1995 ), .C(\U1/keyexpantion/SB0/n1994 ), .D(
        \U1/keyexpantion/SB0/n1993 ), .E(\U1/keyexpantion/SB0/n1992 ), .F(
        \U1/keyexpantion/SB0/n1991 ), .Y(\U1/keyexpantion/ws [13]) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1142  ( .A0(
        \U1/keyexpantion/SB0/n3352 ), .A1(\U1/keyexpantion/SB0/n3305 ), .B0(
        \U1/keyexpantion/SB0/n3310 ), .B1(\U1/keyexpantion/SB0/n2077 ), .C0(
        \U1/keyexpantion/SB0/n1996 ), .Y(\U1/keyexpantion/SB0/n2005 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1141  ( .A0(
        \U1/keyexpantion/SB0/n3284 ), .A1(\U1/keyexpantion/SB0/n2075 ), .B0(
        \U1/keyexpantion/SB0/n3331 ), .Y(\U1/keyexpantion/SB0/n2000 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1140  ( .A0(
        \U1/keyexpantion/SB0/n2062 ), .A1(\U1/keyexpantion/SB0/n3308 ), .B0(
        \U1/keyexpantion/SB0/n2067 ), .Y(\U1/keyexpantion/SB0/n1999 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1139  ( .A(
        \U1/keyexpantion/SB0/n2017 ), .B(\U1/keyexpantion/SB0/n3355 ), .Y(
        \U1/keyexpantion/SB0/n3337 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1138  ( .A0(
        \U1/keyexpantion/SB0/n3314 ), .A1(\U1/keyexpantion/SB0/n3277 ), .B0(
        \U1/keyexpantion/SB0/n3337 ), .Y(\U1/keyexpantion/SB0/n1998 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1137  ( .A(
        \U1/keyexpantion/SB0/n2000 ), .B(\U1/keyexpantion/SB0/n1999 ), .C(
        \U1/keyexpantion/SB0/n1998 ), .D(\U1/keyexpantion/SB0/n1997 ), .Y(
        \U1/keyexpantion/SB0/n2004 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1136  ( .A(
        \U1/keyexpantion/SB0/n3352 ), .B(\U1/keyexpantion/SB0/n3353 ), .Y(
        \U1/keyexpantion/SB0/n2073 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1135  ( .A(
        \U1/keyexpantion/SB0/n3341 ), .B(\U1/keyexpantion/SB0/n2073 ), .Y(
        \U1/keyexpantion/SB0/n2001 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1134  ( .A0(
        \U1/keyexpantion/SB0/n2064 ), .A1(\U1/keyexpantion/SB0/n2002 ), .B0(
        \U1/keyexpantion/SB0/n2001 ), .B1(\U1/keyexpantion/SB0/n2017 ), .C0(
        \U1/keyexpantion/SB0/n2015 ), .C1(\U1/keyexpantion/SB0/n2046 ), .Y(
        \U1/keyexpantion/SB0/n2003 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1133  ( .A(\U1/keyexpantion/SB0/n2008 ), .B(\U1/keyexpantion/SB0/n2007 ), .C(\U1/keyexpantion/SB0/n2006 ), .D(
        \U1/keyexpantion/SB0/n2005 ), .E(\U1/keyexpantion/SB0/n2004 ), .F(
        \U1/keyexpantion/SB0/n2003 ), .Y(\U1/keyexpantion/ws [14]) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1132  ( .A0(
        \U1/keyexpantion/SB0/n2009 ), .A1(\U1/keyexpantion/SB0/n3311 ), .B0(
        \U1/keyexpantion/SB0/n2077 ), .Y(\U1/keyexpantion/SB0/n2021 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U1131  ( .A(
        \U1/keyexpantion/SB0/n2012 ), .B(\U1/keyexpantion/SB0/n2011 ), .C(
        \U1/keyexpantion/SB0/n2010 ), .Y(\U1/keyexpantion/SB0/n2020 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U1130  ( .A(
        \U1/keyexpantion/SB0/n2061 ), .B(\U1/keyexpantion/SB0/n2065 ), .C(
        \U1/keyexpantion/SB0/n3291 ), .Y(\U1/keyexpantion/SB0/n2014 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1129  ( .A0(
        \U1/keyexpantion/SB0/n2016 ), .A1(\U1/keyexpantion/SB0/n2015 ), .B0(
        \U1/keyexpantion/SB0/n2014 ), .B1(\U1/keyexpantion/SB0/n2072 ), .C0(
        \U1/keyexpantion/SB0/n2013 ), .C1(\U1/keyexpantion/SB0/n3289 ), .Y(
        \U1/keyexpantion/SB0/n2019 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1128  ( .A0(
        \U1/keyexpantion/SB0/n3352 ), .A1(\U1/keyexpantion/SB0/n2046 ), .B0(
        \U1/keyexpantion/SB0/n3353 ), .B1(\U1/keyexpantion/SB0/n2017 ), .Y(
        \U1/keyexpantion/SB0/n2018 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1127  ( .A(\U1/keyexpantion/SB0/n2023 ), .B(\U1/keyexpantion/SB0/n2022 ), .C(\U1/keyexpantion/SB0/n2021 ), .D(
        \U1/keyexpantion/SB0/n2020 ), .E(\U1/keyexpantion/SB0/n2019 ), .F(
        \U1/keyexpantion/SB0/n2018 ), .Y(\U1/keyexpantion/SB0/n3361 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1126  ( .A0(
        \U1/keyexpantion/SB0/n3287 ), .A1(\U1/keyexpantion/SB0/n3356 ), .B0(
        \U1/keyexpantion/SB0/n2024 ), .Y(\U1/keyexpantion/SB0/n2040 ) );
  AO22_X0P5M_A12TL \U1/keyexpantion/SB0/U1125  ( .A0(
        \U1/keyexpantion/SB0/n2026 ), .A1(\U1/keyexpantion/SB0/n3278 ), .B0(
        \U1/keyexpantion/SB0/n2025 ), .B1(\U1/keyexpantion/SB0/n3338 ), .Y(
        \U1/keyexpantion/SB0/n2039 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1124  ( .A0(
        \U1/keyexpantion/SB0/n3290 ), .A1(\U1/keyexpantion/SB0/n3353 ), .B0(
        \U1/keyexpantion/SB0/n2028 ), .B1(\U1/keyexpantion/SB0/n2027 ), .C0(
        \U1/keyexpantion/SB0/n2046 ), .C1(\U1/keyexpantion/SB0/n2072 ), .Y(
        \U1/keyexpantion/SB0/n2038 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1123  ( .A(\U1/keyexpantion/SB0/n2032 ), .B(\U1/keyexpantion/SB0/n2031 ), .C(\U1/keyexpantion/SB0/n2030 ), .D(
        \U1/keyexpantion/SB0/n2029 ), .Y(\U1/keyexpantion/SB0/n2037 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1122  ( .AN(
        \U1/keyexpantion/SB0/n2035 ), .B(\U1/keyexpantion/SB0/n2034 ), .C(
        \U1/keyexpantion/SB0/n2033 ), .Y(\U1/keyexpantion/SB0/n2036 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1121  ( .A(\U1/keyexpantion/SB0/n2041 ), .B(\U1/keyexpantion/SB0/n2040 ), .C(\U1/keyexpantion/SB0/n2039 ), .D(
        \U1/keyexpantion/SB0/n2038 ), .E(\U1/keyexpantion/SB0/n2037 ), .F(
        \U1/keyexpantion/SB0/n2036 ), .Y(\U1/keyexpantion/SB0/n3303 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1120  ( .A0(
        \U1/keyexpantion/SB0/n3316 ), .A1(\U1/keyexpantion/SB0/n3336 ), .B0(
        \U1/keyexpantion/SB0/n2061 ), .Y(\U1/keyexpantion/SB0/n2045 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1119  ( .A(
        \U1/keyexpantion/SB0/n2045 ), .B(\U1/keyexpantion/SB0/n2044 ), .C(
        \U1/keyexpantion/SB0/n2043 ), .D(\U1/keyexpantion/SB0/n2042 ), .Y(
        \U1/keyexpantion/SB0/n2058 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1118  ( .A0(
        \U1/keyexpantion/SB0/n3310 ), .A1(\U1/keyexpantion/SB0/n2077 ), .B0(
        \U1/keyexpantion/SB0/n3288 ), .B1(\U1/keyexpantion/SB0/n3289 ), .C0(
        \U1/keyexpantion/SB0/n3318 ), .C1(\U1/keyexpantion/SB0/n2046 ), .Y(
        \U1/keyexpantion/SB0/n2057 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1117  ( .A(
        \U1/keyexpantion/SB0/n2050 ), .B(\U1/keyexpantion/SB0/n2049 ), .C(
        \U1/keyexpantion/SB0/n2048 ), .D(\U1/keyexpantion/SB0/n2047 ), .Y(
        \U1/keyexpantion/SB0/n2056 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U1116  ( .A(
        \U1/keyexpantion/SB0/n2054 ), .B(\U1/keyexpantion/SB0/n2053 ), .C(
        \U1/keyexpantion/SB0/n2052 ), .D(\U1/keyexpantion/SB0/n2051 ), .Y(
        \U1/keyexpantion/SB0/n2055 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1115  ( .A(\U1/keyexpantion/SB0/n2058 ), .B(\U1/keyexpantion/SB0/n2057 ), .C(\U1/keyexpantion/SB0/n2056 ), .D(
        \U1/keyexpantion/SB0/n2055 ), .Y(\U1/keyexpantion/SB0/n2059 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1114  ( .A(\U1/keyexpantion/SB0/n2059 ), .Y(\U1/keyexpantion/SB0/n3294 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1113  ( .A0(
        \U1/keyexpantion/SB0/n2062 ), .A1(\U1/keyexpantion/SB0/n3339 ), .B0(
        \U1/keyexpantion/SB0/n2061 ), .B1(\U1/keyexpantion/SB0/n2060 ), .Y(
        \U1/keyexpantion/SB0/n2063 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U1112  ( .A0(
        \U1/keyexpantion/SB0/n2064 ), .A1(\U1/keyexpantion/SB0/n3318 ), .B0(
        \U1/keyexpantion/SB0/n3294 ), .C0(\U1/keyexpantion/SB0/n2063 ), .Y(
        \U1/keyexpantion/SB0/n2080 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U1111  ( .A1N(
        \U1/keyexpantion/SB0/n2066 ), .A0(\U1/keyexpantion/SB0/n2065 ), .B0(
        \U1/keyexpantion/SB0/n3341 ), .Y(\U1/keyexpantion/SB0/n2070 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1110  ( .A0(
        \U1/keyexpantion/SB0/n3336 ), .A1(\U1/keyexpantion/SB0/n3331 ), .B0(
        \U1/keyexpantion/SB0/n2067 ), .Y(\U1/keyexpantion/SB0/n2069 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1109  ( .AN(
        \U1/keyexpantion/SB0/n2071 ), .B(\U1/keyexpantion/SB0/n2070 ), .C(
        \U1/keyexpantion/SB0/n2069 ), .D(\U1/keyexpantion/SB0/n2068 ), .Y(
        \U1/keyexpantion/SB0/n2079 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1108  ( .A(
        \U1/keyexpantion/SB0/n2072 ), .B(\U1/keyexpantion/SB0/n3352 ), .Y(
        \U1/keyexpantion/SB0/n2074 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1107  ( .A0(
        \U1/keyexpantion/SB0/n2075 ), .A1(\U1/keyexpantion/SB0/n2074 ), .B0(
        \U1/keyexpantion/SB0/n3291 ), .B1(\U1/keyexpantion/SB0/n2073 ), .Y(
        \U1/keyexpantion/SB0/n2076 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1106  ( .A0(
        \U1/keyexpantion/SB0/n3290 ), .A1(\U1/keyexpantion/SB0/n3356 ), .B0(
        \U1/keyexpantion/SB0/n2077 ), .B1(\U1/keyexpantion/SB0/n3351 ), .C0(
        \U1/keyexpantion/SB0/n2076 ), .Y(\U1/keyexpantion/SB0/n2078 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U1105  ( .A(\U1/keyexpantion/SB0/n3361 ), .B(\U1/keyexpantion/SB0/n3303 ), .C(\U1/keyexpantion/SB0/n2081 ), .D(
        \U1/keyexpantion/SB0/n2080 ), .E(\U1/keyexpantion/SB0/n2079 ), .F(
        \U1/keyexpantion/SB0/n2078 ), .Y(\U1/keyexpantion/ws [15]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1104  ( .A(\U1/rkey [15]), .B(
        \U1/rkey [14]), .Y(\U1/keyexpantion/SB0/n2100 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1103  ( .A(\U1/rkey [13]), .B(
        \U1/rkey [12]), .Y(\U1/keyexpantion/SB0/n2091 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1102  ( .A(
        \U1/keyexpantion/SB0/n2100 ), .B(\U1/keyexpantion/SB0/n2091 ), .Y(
        \U1/keyexpantion/SB0/n2165 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1101  ( .A(\U1/rkey [9]), .Y(
        \U1/keyexpantion/SB0/n2085 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1100  ( .A(\U1/rkey [8]), .Y(
        \U1/keyexpantion/SB0/n2082 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1099  ( .A(
        \U1/keyexpantion/SB0/n2085 ), .B(\U1/keyexpantion/SB0/n2082 ), .Y(
        \U1/keyexpantion/SB0/n2092 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1098  ( .A(\U1/rkey [11]), .B(
        \U1/rkey [10]), .Y(\U1/keyexpantion/SB0/n2112 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1097  ( .A(
        \U1/keyexpantion/SB0/n2092 ), .B(\U1/keyexpantion/SB0/n2112 ), .Y(
        \U1/keyexpantion/SB0/n2472 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1096  ( .A(
        \U1/keyexpantion/SB0/n2165 ), .B(\U1/keyexpantion/SB0/n2472 ), .Y(
        \U1/keyexpantion/SB0/n2254 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U1095  ( .A(\U1/rkey [10]), .B(
        \U1/rkey [11]), .Y(\U1/keyexpantion/SB0/n2095 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1094  ( .A(
        \U1/keyexpantion/SB0/n2095 ), .B(\U1/keyexpantion/SB0/n2092 ), .Y(
        \U1/keyexpantion/SB0/n2410 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1093  ( .A(\U1/rkey [15]), .Y(
        \U1/keyexpantion/SB0/n2088 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1092  ( .A(
        \U1/keyexpantion/SB0/n2088 ), .B(\U1/rkey [14]), .Y(
        \U1/keyexpantion/SB0/n2118 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1091  ( .A(
        \U1/keyexpantion/SB0/n2118 ), .B(\U1/keyexpantion/SB0/n2091 ), .Y(
        \U1/keyexpantion/SB0/n2164 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1090  ( .A(
        \U1/keyexpantion/SB0/n2410 ), .B(\U1/keyexpantion/SB0/n2164 ), .Y(
        \U1/keyexpantion/SB0/n2376 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1089  ( .A(\U1/rkey [11]), .Y(
        \U1/keyexpantion/SB0/n2083 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U1088  ( .A(\U1/rkey [10]), .B(
        \U1/keyexpantion/SB0/n2083 ), .Y(\U1/keyexpantion/SB0/n2093 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1087  ( .A(
        \U1/keyexpantion/SB0/n2092 ), .B(\U1/keyexpantion/SB0/n2093 ), .Y(
        \U1/keyexpantion/SB0/n2316 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1086  ( .A(\U1/keyexpantion/SB0/n2316 ), .Y(\U1/keyexpantion/SB0/n2506 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1085  ( .A(\U1/rkey [12]), .Y(
        \U1/keyexpantion/SB0/n2084 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1084  ( .A(
        \U1/keyexpantion/SB0/n2084 ), .B(\U1/rkey [13]), .Y(
        \U1/keyexpantion/SB0/n2099 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1083  ( .A(\U1/rkey [14]), .Y(
        \U1/keyexpantion/SB0/n2087 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1082  ( .A(
        \U1/keyexpantion/SB0/n2087 ), .B(\U1/rkey [15]), .Y(
        \U1/keyexpantion/SB0/n2109 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1081  ( .A(
        \U1/keyexpantion/SB0/n2099 ), .B(\U1/keyexpantion/SB0/n2109 ), .Y(
        \U1/keyexpantion/SB0/n2362 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1080  ( .A(\U1/keyexpantion/SB0/n2362 ), .Y(\U1/keyexpantion/SB0/n2460 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1079  ( .A(
        \U1/keyexpantion/SB0/n2506 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2294 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1078  ( .A(\U1/keyexpantion/SB0/n2165 ), .Y(\U1/keyexpantion/SB0/n2475 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1077  ( .A(\U1/rkey [9]), .B(
        \U1/rkey [8]), .Y(\U1/keyexpantion/SB0/n2096 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1076  ( .A(
        \U1/keyexpantion/SB0/n2096 ), .B(\U1/keyexpantion/SB0/n2112 ), .Y(
        \U1/keyexpantion/SB0/n2428 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1075  ( .A(\U1/keyexpantion/SB0/n2428 ), .Y(\U1/keyexpantion/SB0/n2516 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1074  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2516 ), .Y(
        \U1/keyexpantion/SB0/n2433 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1073  ( .A(
        \U1/keyexpantion/SB0/n2082 ), .B(\U1/rkey [9]), .Y(
        \U1/keyexpantion/SB0/n2111 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1072  ( .A(
        \U1/keyexpantion/SB0/n2093 ), .B(\U1/keyexpantion/SB0/n2111 ), .Y(
        \U1/keyexpantion/SB0/n2303 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1071  ( .A(\U1/keyexpantion/SB0/n2303 ), .Y(\U1/keyexpantion/SB0/n2417 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1070  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2272 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U1069  ( .A(
        \U1/keyexpantion/SB0/n2294 ), .B(\U1/keyexpantion/SB0/n2433 ), .C(
        \U1/keyexpantion/SB0/n2272 ), .Y(\U1/keyexpantion/SB0/n2131 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1068  ( .A(
        \U1/keyexpantion/SB0/n2091 ), .B(\U1/keyexpantion/SB0/n2109 ), .Y(
        \U1/keyexpantion/SB0/n2361 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1067  ( .A(
        \U1/keyexpantion/SB0/n2083 ), .B(\U1/rkey [10]), .Y(
        \U1/keyexpantion/SB0/n2102 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1066  ( .A(
        \U1/keyexpantion/SB0/n2102 ), .B(\U1/keyexpantion/SB0/n2111 ), .Y(
        \U1/keyexpantion/SB0/n2359 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1065  ( .A(
        \U1/keyexpantion/SB0/n2361 ), .B(\U1/keyexpantion/SB0/n2359 ), .Y(
        \U1/keyexpantion/SB0/n2249 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1064  ( .A(\U1/keyexpantion/SB0/n2164 ), .Y(\U1/keyexpantion/SB0/n2477 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1063  ( .A(\U1/rkey [13]), .Y(
        \U1/keyexpantion/SB0/n2086 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1062  ( .A(
        \U1/keyexpantion/SB0/n2084 ), .B(\U1/keyexpantion/SB0/n2086 ), .Y(
        \U1/keyexpantion/SB0/n2110 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1061  ( .A(
        \U1/keyexpantion/SB0/n2100 ), .B(\U1/keyexpantion/SB0/n2110 ), .Y(
        \U1/keyexpantion/SB0/n2520 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1060  ( .A(\U1/keyexpantion/SB0/n2520 ), .Y(\U1/keyexpantion/SB0/n2451 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1059  ( .A(
        \U1/keyexpantion/SB0/n2085 ), .B(\U1/rkey [8]), .Y(
        \U1/keyexpantion/SB0/n2101 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1058  ( .A(
        \U1/keyexpantion/SB0/n2101 ), .B(\U1/keyexpantion/SB0/n2112 ), .Y(
        \U1/keyexpantion/SB0/n2485 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1057  ( .A(\U1/keyexpantion/SB0/n2485 ), .Y(\U1/keyexpantion/SB0/n2308 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1056  ( .A0(
        \U1/keyexpantion/SB0/n2477 ), .A1(\U1/keyexpantion/SB0/n2451 ), .B0(
        \U1/keyexpantion/SB0/n2308 ), .Y(\U1/keyexpantion/SB0/n2090 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1055  ( .A(
        \U1/keyexpantion/SB0/n2096 ), .B(\U1/keyexpantion/SB0/n2093 ), .Y(
        \U1/keyexpantion/SB0/n2473 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1054  ( .A(\U1/keyexpantion/SB0/n2473 ), .Y(\U1/keyexpantion/SB0/n2459 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1053  ( .A(
        \U1/keyexpantion/SB0/n2086 ), .B(\U1/rkey [12]), .Y(
        \U1/keyexpantion/SB0/n2117 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1052  ( .A(
        \U1/keyexpantion/SB0/n2109 ), .B(\U1/keyexpantion/SB0/n2117 ), .Y(
        \U1/keyexpantion/SB0/n2513 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1051  ( .A(
        \U1/keyexpantion/SB0/n2361 ), .B(\U1/keyexpantion/SB0/n2513 ), .Y(
        \U1/keyexpantion/SB0/n2227 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1050  ( .A(
        \U1/keyexpantion/SB0/n2088 ), .B(\U1/keyexpantion/SB0/n2087 ), .Y(
        \U1/keyexpantion/SB0/n2108 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1049  ( .A(
        \U1/keyexpantion/SB0/n2099 ), .B(\U1/keyexpantion/SB0/n2108 ), .Y(
        \U1/keyexpantion/SB0/n2488 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1048  ( .A(\U1/keyexpantion/SB0/n2488 ), .Y(\U1/keyexpantion/SB0/n2208 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1047  ( .A0(
        \U1/keyexpantion/SB0/n2459 ), .A1(\U1/keyexpantion/SB0/n2227 ), .B0(
        \U1/keyexpantion/SB0/n2208 ), .B1(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2089 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U1046  ( .AN(
        \U1/keyexpantion/SB0/n2249 ), .B(\U1/keyexpantion/SB0/n2090 ), .C(
        \U1/keyexpantion/SB0/n2089 ), .Y(\U1/keyexpantion/SB0/n2130 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1045  ( .A(
        \U1/keyexpantion/SB0/n2091 ), .B(\U1/keyexpantion/SB0/n2108 ), .Y(
        \U1/keyexpantion/SB0/n2378 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1044  ( .A(
        \U1/keyexpantion/SB0/n2095 ), .B(\U1/keyexpantion/SB0/n2096 ), .Y(
        \U1/keyexpantion/SB0/n2523 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1043  ( .A(
        \U1/keyexpantion/SB0/n2118 ), .B(\U1/keyexpantion/SB0/n2099 ), .Y(
        \U1/keyexpantion/SB0/n2429 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1042  ( .A(
        \U1/keyexpantion/SB0/n2095 ), .B(\U1/keyexpantion/SB0/n2101 ), .Y(
        \U1/keyexpantion/SB0/n2426 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1041  ( .A(
        \U1/keyexpantion/SB0/n2092 ), .B(\U1/keyexpantion/SB0/n2102 ), .Y(
        \U1/keyexpantion/SB0/n2431 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1040  ( .A(\U1/keyexpantion/SB0/n2431 ), .Y(\U1/keyexpantion/SB0/n2411 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1039  ( .A(\U1/keyexpantion/SB0/n2513 ), .Y(\U1/keyexpantion/SB0/n2222 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1038  ( .A(
        \U1/keyexpantion/SB0/n2093 ), .B(\U1/keyexpantion/SB0/n2101 ), .Y(
        \U1/keyexpantion/SB0/n2449 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1037  ( .A(\U1/keyexpantion/SB0/n2449 ), .Y(\U1/keyexpantion/SB0/n2474 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U1036  ( .A0(
        \U1/keyexpantion/SB0/n2411 ), .A1(\U1/keyexpantion/SB0/n2475 ), .B0(
        \U1/keyexpantion/SB0/n2222 ), .B1(\U1/keyexpantion/SB0/n2474 ), .Y(
        \U1/keyexpantion/SB0/n2094 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U1035  ( .A0(
        \U1/keyexpantion/SB0/n2378 ), .A1(\U1/keyexpantion/SB0/n2523 ), .B0(
        \U1/keyexpantion/SB0/n2429 ), .B1(\U1/keyexpantion/SB0/n2426 ), .C0(
        \U1/keyexpantion/SB0/n2094 ), .Y(\U1/keyexpantion/SB0/n2129 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1034  ( .A(
        \U1/keyexpantion/SB0/n2431 ), .B(\U1/keyexpantion/SB0/n2378 ), .Y(
        \U1/keyexpantion/SB0/n2215 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1033  ( .A(
        \U1/keyexpantion/SB0/n2426 ), .B(\U1/keyexpantion/SB0/n2361 ), .Y(
        \U1/keyexpantion/SB0/n2225 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1032  ( .A(\U1/keyexpantion/SB0/n2225 ), .Y(\U1/keyexpantion/SB0/n2098 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1031  ( .A(
        \U1/keyexpantion/SB0/n2095 ), .B(\U1/keyexpantion/SB0/n2111 ), .Y(
        \U1/keyexpantion/SB0/n2501 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1030  ( .A(\U1/keyexpantion/SB0/n2501 ), .Y(\U1/keyexpantion/SB0/n2450 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1029  ( .A(
        \U1/keyexpantion/SB0/n2096 ), .B(\U1/keyexpantion/SB0/n2102 ), .Y(
        \U1/keyexpantion/SB0/n2486 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1028  ( .A(\U1/keyexpantion/SB0/n2486 ), .Y(\U1/keyexpantion/SB0/n2497 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U1027  ( .A0(
        \U1/keyexpantion/SB0/n2450 ), .A1(\U1/keyexpantion/SB0/n2497 ), .B0(
        \U1/keyexpantion/SB0/n2451 ), .Y(\U1/keyexpantion/SB0/n2097 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1026  ( .A(
        \U1/keyexpantion/SB0/n2100 ), .B(\U1/keyexpantion/SB0/n2117 ), .Y(
        \U1/keyexpantion/SB0/n2502 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1025  ( .A(\U1/keyexpantion/SB0/n2502 ), .Y(\U1/keyexpantion/SB0/n2452 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1024  ( .A(
        \U1/keyexpantion/SB0/n2452 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2242 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1023  ( .AN(
        \U1/keyexpantion/SB0/n2215 ), .B(\U1/keyexpantion/SB0/n2098 ), .C(
        \U1/keyexpantion/SB0/n2097 ), .D(\U1/keyexpantion/SB0/n2242 ), .Y(
        \U1/keyexpantion/SB0/n2107 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1022  ( .A(
        \U1/keyexpantion/SB0/n2110 ), .B(\U1/keyexpantion/SB0/n2108 ), .Y(
        \U1/keyexpantion/SB0/n2522 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1021  ( .A(
        \U1/keyexpantion/SB0/n2100 ), .B(\U1/keyexpantion/SB0/n2099 ), .Y(
        \U1/keyexpantion/SB0/n2514 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U1020  ( .A0(
        \U1/keyexpantion/SB0/n2164 ), .A1(\U1/keyexpantion/SB0/n2316 ), .B0(
        \U1/keyexpantion/SB0/n2522 ), .B1(\U1/keyexpantion/SB0/n2431 ), .C0(
        \U1/keyexpantion/SB0/n2514 ), .C1(\U1/keyexpantion/SB0/n2449 ), .Y(
        \U1/keyexpantion/SB0/n2106 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1019  ( .A(
        \U1/keyexpantion/SB0/n2473 ), .B(\U1/keyexpantion/SB0/n2164 ), .Y(
        \U1/keyexpantion/SB0/n2300 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1018  ( .A(
        \U1/keyexpantion/SB0/n2222 ), .B(\U1/keyexpantion/SB0/n2411 ), .Y(
        \U1/keyexpantion/SB0/n2253 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1017  ( .A(
        \U1/keyexpantion/SB0/n2474 ), .B(\U1/keyexpantion/SB0/n2475 ), .Y(
        \U1/keyexpantion/SB0/n2273 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1016  ( .A(\U1/keyexpantion/SB0/n2429 ), .Y(\U1/keyexpantion/SB0/n2503 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1015  ( .A(
        \U1/keyexpantion/SB0/n2503 ), .B(\U1/keyexpantion/SB0/n2308 ), .Y(
        \U1/keyexpantion/SB0/n2311 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1014  ( .AN(
        \U1/keyexpantion/SB0/n2300 ), .B(\U1/keyexpantion/SB0/n2253 ), .C(
        \U1/keyexpantion/SB0/n2273 ), .D(\U1/keyexpantion/SB0/n2311 ), .Y(
        \U1/keyexpantion/SB0/n2105 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1013  ( .A(
        \U1/keyexpantion/SB0/n2118 ), .B(\U1/keyexpantion/SB0/n2110 ), .Y(
        \U1/keyexpantion/SB0/n2223 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1012  ( .A(
        \U1/keyexpantion/SB0/n2223 ), .B(\U1/keyexpantion/SB0/n2485 ), .Y(
        \U1/keyexpantion/SB0/n2402 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1011  ( .A(
        \U1/keyexpantion/SB0/n2102 ), .B(\U1/keyexpantion/SB0/n2101 ), .Y(
        \U1/keyexpantion/SB0/n2521 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1010  ( .A(
        \U1/keyexpantion/SB0/n2488 ), .B(\U1/keyexpantion/SB0/n2521 ), .Y(
        \U1/keyexpantion/SB0/n2367 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1009  ( .A(\U1/keyexpantion/SB0/n2367 ), .Y(\U1/keyexpantion/SB0/n2103 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1008  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2308 ), .Y(
        \U1/keyexpantion/SB0/n2386 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1007  ( .A(\U1/keyexpantion/SB0/n2521 ), .Y(\U1/keyexpantion/SB0/n2504 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1006  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2504 ), .Y(
        \U1/keyexpantion/SB0/n2437 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U1005  ( .AN(
        \U1/keyexpantion/SB0/n2402 ), .B(\U1/keyexpantion/SB0/n2103 ), .C(
        \U1/keyexpantion/SB0/n2386 ), .D(\U1/keyexpantion/SB0/n2437 ), .Y(
        \U1/keyexpantion/SB0/n2104 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U1004  ( .A(\U1/keyexpantion/SB0/n2107 ), .B(\U1/keyexpantion/SB0/n2106 ), .C(\U1/keyexpantion/SB0/n2105 ), .D(
        \U1/keyexpantion/SB0/n2104 ), .Y(\U1/keyexpantion/SB0/n2204 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1003  ( .A(
        \U1/keyexpantion/SB0/n2428 ), .B(\U1/keyexpantion/SB0/n2223 ), .Y(
        \U1/keyexpantion/SB0/n2436 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U1002  ( .A(
        \U1/keyexpantion/SB0/n2117 ), .B(\U1/keyexpantion/SB0/n2108 ), .Y(
        \U1/keyexpantion/SB0/n2319 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U1001  ( .A(
        \U1/keyexpantion/SB0/n2410 ), .B(\U1/keyexpantion/SB0/n2319 ), .Y(
        \U1/keyexpantion/SB0/n2290 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U1000  ( .A(\U1/keyexpantion/SB0/n2522 ), .Y(\U1/keyexpantion/SB0/n2478 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U999  ( .A(
        \U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2459 ), .Y(
        \U1/keyexpantion/SB0/n2239 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U998  ( .A0(
        \U1/keyexpantion/SB0/n2319 ), .A1(\U1/keyexpantion/SB0/n2521 ), .B0(
        \U1/keyexpantion/SB0/n2239 ), .Y(\U1/keyexpantion/SB0/n2116 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U997  ( .A(\U1/keyexpantion/SB0/n2359 ), 
        .Y(\U1/keyexpantion/SB0/n2454 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U996  ( .A(
        \U1/keyexpantion/SB0/n2454 ), .B(\U1/keyexpantion/SB0/n2477 ), .Y(
        \U1/keyexpantion/SB0/n2455 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U995  ( .A(
        \U1/keyexpantion/SB0/n2477 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2414 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U994  ( .A(
        \U1/keyexpantion/SB0/n2110 ), .B(\U1/keyexpantion/SB0/n2109 ), .Y(
        \U1/keyexpantion/SB0/n2484 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U993  ( .A(\U1/keyexpantion/SB0/n2484 ), 
        .Y(\U1/keyexpantion/SB0/n2234 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U992  ( .A(
        \U1/keyexpantion/SB0/n2450 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2258 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U991  ( .A(\U1/keyexpantion/SB0/n2472 ), 
        .Y(\U1/keyexpantion/SB0/n2453 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U990  ( .A(
        \U1/keyexpantion/SB0/n2453 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2322 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U989  ( .A(
        \U1/keyexpantion/SB0/n2455 ), .B(\U1/keyexpantion/SB0/n2414 ), .C(
        \U1/keyexpantion/SB0/n2258 ), .D(\U1/keyexpantion/SB0/n2322 ), .Y(
        \U1/keyexpantion/SB0/n2115 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U988  ( .A(
        \U1/keyexpantion/SB0/n2474 ), .B(\U1/keyexpantion/SB0/n2452 ), .Y(
        \U1/keyexpantion/SB0/n2381 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U987  ( .A(
        \U1/keyexpantion/SB0/n2516 ), .B(\U1/keyexpantion/SB0/n2452 ), .Y(
        \U1/keyexpantion/SB0/n2372 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U986  ( .A(\U1/keyexpantion/SB0/n2514 ), 
        .Y(\U1/keyexpantion/SB0/n2507 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U985  ( .A(
        \U1/keyexpantion/SB0/n2411 ), .B(\U1/keyexpantion/SB0/n2507 ), .Y(
        \U1/keyexpantion/SB0/n2219 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U984  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2450 ), .Y(
        \U1/keyexpantion/SB0/n2355 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U983  ( .A(
        \U1/keyexpantion/SB0/n2381 ), .B(\U1/keyexpantion/SB0/n2372 ), .C(
        \U1/keyexpantion/SB0/n2219 ), .D(\U1/keyexpantion/SB0/n2355 ), .Y(
        \U1/keyexpantion/SB0/n2114 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U982  ( .A(\U1/keyexpantion/SB0/n2426 ), 
        .Y(\U1/keyexpantion/SB0/n2395 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U981  ( .A(
        \U1/keyexpantion/SB0/n2222 ), .B(\U1/keyexpantion/SB0/n2395 ), .Y(
        \U1/keyexpantion/SB0/n2206 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U980  ( .A(
        \U1/keyexpantion/SB0/n2112 ), .B(\U1/keyexpantion/SB0/n2111 ), .Y(
        \U1/keyexpantion/SB0/n2461 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U979  ( .A(\U1/keyexpantion/SB0/n2461 ), 
        .Y(\U1/keyexpantion/SB0/n2495 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U978  ( .A(
        \U1/keyexpantion/SB0/n2222 ), .B(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2270 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U977  ( .A(\U1/keyexpantion/SB0/n2410 ), 
        .Y(\U1/keyexpantion/SB0/n2518 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U976  ( .A(
        \U1/keyexpantion/SB0/n2518 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2305 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U975  ( .A(
        \U1/keyexpantion/SB0/n2451 ), .B(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2479 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U974  ( .A(
        \U1/keyexpantion/SB0/n2206 ), .B(\U1/keyexpantion/SB0/n2270 ), .C(
        \U1/keyexpantion/SB0/n2305 ), .D(\U1/keyexpantion/SB0/n2479 ), .Y(
        \U1/keyexpantion/SB0/n2113 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U973  ( .A(\U1/keyexpantion/SB0/n2436 ), 
        .B(\U1/keyexpantion/SB0/n2290 ), .C(\U1/keyexpantion/SB0/n2116 ), .D(
        \U1/keyexpantion/SB0/n2115 ), .E(\U1/keyexpantion/SB0/n2114 ), .F(
        \U1/keyexpantion/SB0/n2113 ), .Y(\U1/keyexpantion/SB0/n2193 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U972  ( .A(\U1/keyexpantion/SB0/n2193 ), 
        .Y(\U1/keyexpantion/SB0/n2127 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U971  ( .A(\U1/keyexpantion/SB0/n2486 ), .B(\U1/keyexpantion/SB0/n2319 ), .Y(\U1/keyexpantion/SB0/n2216 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U970  ( .A(
        \U1/keyexpantion/SB0/n2118 ), .B(\U1/keyexpantion/SB0/n2117 ), .Y(
        \U1/keyexpantion/SB0/n2483 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U969  ( .A(\U1/keyexpantion/SB0/n2483 ), .B(\U1/keyexpantion/SB0/n2359 ), .Y(\U1/keyexpantion/SB0/n2368 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U968  ( .A(\U1/keyexpantion/SB0/n2368 ), 
        .Y(\U1/keyexpantion/SB0/n2120 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U967  ( .A(\U1/keyexpantion/SB0/n2361 ), 
        .Y(\U1/keyexpantion/SB0/n2508 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U966  ( .A0(
        \U1/keyexpantion/SB0/n2234 ), .A1(\U1/keyexpantion/SB0/n2508 ), .B0(
        \U1/keyexpantion/SB0/n2495 ), .Y(\U1/keyexpantion/SB0/n2119 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U965  ( .A(
        \U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2395 ), .Y(
        \U1/keyexpantion/SB0/n2241 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U964  ( .AN(
        \U1/keyexpantion/SB0/n2216 ), .B(\U1/keyexpantion/SB0/n2120 ), .C(
        \U1/keyexpantion/SB0/n2119 ), .D(\U1/keyexpantion/SB0/n2241 ), .Y(
        \U1/keyexpantion/SB0/n2124 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U963  ( .A0(
        \U1/keyexpantion/SB0/n2472 ), .A1(\U1/keyexpantion/SB0/n2520 ), .B0(
        \U1/keyexpantion/SB0/n2378 ), .B1(\U1/keyexpantion/SB0/n2426 ), .C0(
        \U1/keyexpantion/SB0/n2485 ), .C1(\U1/keyexpantion/SB0/n2502 ), .Y(
        \U1/keyexpantion/SB0/n2123 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U962  ( .A(\U1/keyexpantion/SB0/n2520 ), .B(\U1/keyexpantion/SB0/n2523 ), .Y(\U1/keyexpantion/SB0/n2281 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U961  ( .A(
        \U1/keyexpantion/SB0/n2508 ), .B(\U1/keyexpantion/SB0/n2450 ), .Y(
        \U1/keyexpantion/SB0/n2439 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U960  ( .A(
        \U1/keyexpantion/SB0/n2411 ), .B(\U1/keyexpantion/SB0/n2508 ), .Y(
        \U1/keyexpantion/SB0/n2373 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U959  ( .A(
        \U1/keyexpantion/SB0/n2395 ), .B(\U1/keyexpantion/SB0/n2475 ), .Y(
        \U1/keyexpantion/SB0/n2220 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U958  ( .AN(
        \U1/keyexpantion/SB0/n2281 ), .B(\U1/keyexpantion/SB0/n2439 ), .C(
        \U1/keyexpantion/SB0/n2373 ), .D(\U1/keyexpantion/SB0/n2220 ), .Y(
        \U1/keyexpantion/SB0/n2122 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U957  ( .A(
        \U1/keyexpantion/SB0/n2518 ), .B(\U1/keyexpantion/SB0/n2503 ), .Y(
        \U1/keyexpantion/SB0/n2293 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U956  ( .A(
        \U1/keyexpantion/SB0/n2395 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2385 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U955  ( .A(
        \U1/keyexpantion/SB0/n2222 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2261 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U954  ( .A(
        \U1/keyexpantion/SB0/n2454 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2306 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U953  ( .A(
        \U1/keyexpantion/SB0/n2293 ), .B(\U1/keyexpantion/SB0/n2385 ), .C(
        \U1/keyexpantion/SB0/n2261 ), .D(\U1/keyexpantion/SB0/n2306 ), .Y(
        \U1/keyexpantion/SB0/n2121 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U952  ( .A(\U1/keyexpantion/SB0/n2124 ), 
        .B(\U1/keyexpantion/SB0/n2123 ), .C(\U1/keyexpantion/SB0/n2122 ), .D(
        \U1/keyexpantion/SB0/n2121 ), .Y(\U1/keyexpantion/SB0/n2125 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U951  ( .A(\U1/keyexpantion/SB0/n2125 ), 
        .Y(\U1/keyexpantion/SB0/n2500 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U950  ( .A(
        \U1/keyexpantion/SB0/n2516 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2126 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U949  ( .AN(
        \U1/keyexpantion/SB0/n2204 ), .B(\U1/keyexpantion/SB0/n2127 ), .C(
        \U1/keyexpantion/SB0/n2500 ), .D(\U1/keyexpantion/SB0/n2126 ), .Y(
        \U1/keyexpantion/SB0/n2128 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U948  ( .A(\U1/keyexpantion/SB0/n2254 ), 
        .B(\U1/keyexpantion/SB0/n2376 ), .C(\U1/keyexpantion/SB0/n2131 ), .D(
        \U1/keyexpantion/SB0/n2130 ), .E(\U1/keyexpantion/SB0/n2129 ), .F(
        \U1/keyexpantion/SB0/n2128 ), .Y(\U1/keyexpantion/SB0/n2183 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U947  ( .A(\U1/keyexpantion/SB0/n2501 ), .B(\U1/keyexpantion/SB0/n2164 ), .Y(\U1/keyexpantion/SB0/n2299 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U946  ( .A(
        \U1/keyexpantion/SB0/n2451 ), .B(\U1/keyexpantion/SB0/n2518 ), .Y(
        \U1/keyexpantion/SB0/n2375 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U945  ( .A(
        \U1/keyexpantion/SB0/n2507 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2252 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U944  ( .A(\U1/keyexpantion/SB0/n2223 ), 
        .Y(\U1/keyexpantion/SB0/n2496 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U943  ( .A(
        \U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2275 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U942  ( .AN(
        \U1/keyexpantion/SB0/n2299 ), .B(\U1/keyexpantion/SB0/n2375 ), .C(
        \U1/keyexpantion/SB0/n2252 ), .D(\U1/keyexpantion/SB0/n2275 ), .Y(
        \U1/keyexpantion/SB0/n2138 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U941  ( .A(\U1/keyexpantion/SB0/n2488 ), .B(\U1/keyexpantion/SB0/n2359 ), .Y(\U1/keyexpantion/SB0/n2401 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U940  ( .A(
        \U1/keyexpantion/SB0/n2411 ), .B(\U1/keyexpantion/SB0/n2477 ), .Y(
        \U1/keyexpantion/SB0/n2232 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U939  ( .A0(
        \U1/keyexpantion/SB0/n2497 ), .A1(\U1/keyexpantion/SB0/n2417 ), .B0(
        \U1/keyexpantion/SB0/n2222 ), .Y(\U1/keyexpantion/SB0/n2132 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U938  ( .A(
        \U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2324 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U937  ( .AN(
        \U1/keyexpantion/SB0/n2401 ), .B(\U1/keyexpantion/SB0/n2232 ), .C(
        \U1/keyexpantion/SB0/n2132 ), .D(\U1/keyexpantion/SB0/n2324 ), .Y(
        \U1/keyexpantion/SB0/n2133 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U936  ( .A(\U1/keyexpantion/SB0/n2133 ), 
        .Y(\U1/keyexpantion/SB0/n2137 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U935  ( .A(\U1/keyexpantion/SB0/n2378 ), 
        .Y(\U1/keyexpantion/SB0/n2498 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U934  ( .A(\U1/keyexpantion/SB0/n2523 ), 
        .Y(\U1/keyexpantion/SB0/n2418 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U933  ( .A0(
        \U1/keyexpantion/SB0/n2518 ), .A1(\U1/keyexpantion/SB0/n2452 ), .B0(
        \U1/keyexpantion/SB0/n2498 ), .B1(\U1/keyexpantion/SB0/n2308 ), .C0(
        \U1/keyexpantion/SB0/n2418 ), .C1(\U1/keyexpantion/SB0/n2496 ), .Y(
        \U1/keyexpantion/SB0/n2136 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U932  ( .A0(
        \U1/keyexpantion/SB0/n2319 ), .A1(\U1/keyexpantion/SB0/n2501 ), .B0(
        \U1/keyexpantion/SB0/n2521 ), .B1(\U1/keyexpantion/SB0/n2522 ), .Y(
        \U1/keyexpantion/SB0/n2134 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U931  ( .A0(
        \U1/keyexpantion/SB0/n2395 ), .A1(\U1/keyexpantion/SB0/n2208 ), .B0(
        \U1/keyexpantion/SB0/n2451 ), .B1(\U1/keyexpantion/SB0/n2474 ), .C0(
        \U1/keyexpantion/SB0/n2134 ), .Y(\U1/keyexpantion/SB0/n2135 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U930  ( .AN(
        \U1/keyexpantion/SB0/n2138 ), .B(\U1/keyexpantion/SB0/n2137 ), .C(
        \U1/keyexpantion/SB0/n2136 ), .D(\U1/keyexpantion/SB0/n2135 ), .Y(
        \U1/keyexpantion/SB0/n2202 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U929  ( .A(\U1/keyexpantion/SB0/n2522 ), .B(\U1/keyexpantion/SB0/n2359 ), .Y(\U1/keyexpantion/SB0/n2217 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U928  ( .A0(
        \U1/keyexpantion/SB0/n2429 ), .A1(\U1/keyexpantion/SB0/n2522 ), .B0(
        \U1/keyexpantion/SB0/n2461 ), .Y(\U1/keyexpantion/SB0/n2143 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U927  ( .A(
        \U1/keyexpantion/SB0/n2461 ), .B(\U1/keyexpantion/SB0/n2449 ), .Y(
        \U1/keyexpantion/SB0/n2301 ) );
  AO22_X0P5M_A12TL \U1/keyexpantion/SB0/U926  ( .A0(
        \U1/keyexpantion/SB0/n2450 ), .A1(\U1/keyexpantion/SB0/n2208 ), .B0(
        \U1/keyexpantion/SB0/n2301 ), .B1(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2142 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U925  ( .A0(
        \U1/keyexpantion/SB0/n2483 ), .A1(\U1/keyexpantion/SB0/n2523 ), .B0(
        \U1/keyexpantion/SB0/n2223 ), .B1(\U1/keyexpantion/SB0/n2316 ), .C0(
        \U1/keyexpantion/SB0/n2485 ), .C1(\U1/keyexpantion/SB0/n2514 ), .Y(
        \U1/keyexpantion/SB0/n2141 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U924  ( .A(\U1/keyexpantion/SB0/n2319 ), 
        .Y(\U1/keyexpantion/SB0/n2412 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U923  ( .A(
        \U1/keyexpantion/SB0/n2516 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2438 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U922  ( .A(
        \U1/keyexpantion/SB0/n2411 ), .B(\U1/keyexpantion/SB0/n2208 ), .Y(
        \U1/keyexpantion/SB0/n2240 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U921  ( .A(
        \U1/keyexpantion/SB0/n2222 ), .B(\U1/keyexpantion/SB0/n2454 ), .Y(
        \U1/keyexpantion/SB0/n2260 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U920  ( .A(
        \U1/keyexpantion/SB0/n2411 ), .B(\U1/keyexpantion/SB0/n2452 ), .Y(
        \U1/keyexpantion/SB0/n2384 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U919  ( .A(
        \U1/keyexpantion/SB0/n2438 ), .B(\U1/keyexpantion/SB0/n2240 ), .C(
        \U1/keyexpantion/SB0/n2260 ), .D(\U1/keyexpantion/SB0/n2384 ), .Y(
        \U1/keyexpantion/SB0/n2140 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U918  ( .A(\U1/keyexpantion/SB0/n2431 ), .B(\U1/keyexpantion/SB0/n2319 ), .Y(\U1/keyexpantion/SB0/n2282 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U917  ( .A(
        \U1/keyexpantion/SB0/n2417 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2292 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U916  ( .A(
        \U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2308 ), .Y(
        \U1/keyexpantion/SB0/n2323 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U915  ( .AN(
        \U1/keyexpantion/SB0/n2282 ), .B(\U1/keyexpantion/SB0/n2292 ), .C(
        \U1/keyexpantion/SB0/n2323 ), .Y(\U1/keyexpantion/SB0/n2139 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U914  ( .A(\U1/keyexpantion/SB0/n2217 ), 
        .B(\U1/keyexpantion/SB0/n2143 ), .C(\U1/keyexpantion/SB0/n2142 ), .D(
        \U1/keyexpantion/SB0/n2141 ), .E(\U1/keyexpantion/SB0/n2140 ), .F(
        \U1/keyexpantion/SB0/n2139 ), .Y(\U1/keyexpantion/SB0/n2529 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U913  ( .A0(
        \U1/keyexpantion/SB0/n2222 ), .A1(\U1/keyexpantion/SB0/n2475 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2144 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U912  ( .A(
        \U1/keyexpantion/SB0/n2208 ), .B(\U1/keyexpantion/SB0/n2308 ), .Y(
        \U1/keyexpantion/SB0/n2370 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U911  ( .A(
        \U1/keyexpantion/SB0/n2450 ), .B(\U1/keyexpantion/SB0/n2498 ), .Y(
        \U1/keyexpantion/SB0/n2237 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U910  ( .A(
        \U1/keyexpantion/SB0/n2498 ), .B(\U1/keyexpantion/SB0/n2454 ), .Y(
        \U1/keyexpantion/SB0/n2288 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U909  ( .A(
        \U1/keyexpantion/SB0/n2144 ), .B(\U1/keyexpantion/SB0/n2370 ), .C(
        \U1/keyexpantion/SB0/n2237 ), .D(\U1/keyexpantion/SB0/n2288 ), .Y(
        \U1/keyexpantion/SB0/n2148 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U908  ( .A0(
        \U1/keyexpantion/SB0/n2501 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2223 ), .B1(\U1/keyexpantion/SB0/n2473 ), .C0(
        \U1/keyexpantion/SB0/n2502 ), .C1(\U1/keyexpantion/SB0/n2359 ), .Y(
        \U1/keyexpantion/SB0/n2147 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U907  ( .A(
        \U1/keyexpantion/SB0/n2453 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2269 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U906  ( .A(
        \U1/keyexpantion/SB0/n2452 ), .B(\U1/keyexpantion/SB0/n2504 ), .Y(
        \U1/keyexpantion/SB0/n2434 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U905  ( .A(
        \U1/keyexpantion/SB0/n2452 ), .B(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2256 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U904  ( .A(
        \U1/keyexpantion/SB0/n2507 ), .B(\U1/keyexpantion/SB0/n2497 ), .Y(
        \U1/keyexpantion/SB0/n2218 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U903  ( .A(
        \U1/keyexpantion/SB0/n2269 ), .B(\U1/keyexpantion/SB0/n2434 ), .C(
        \U1/keyexpantion/SB0/n2256 ), .D(\U1/keyexpantion/SB0/n2218 ), .Y(
        \U1/keyexpantion/SB0/n2146 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U902  ( .A(
        \U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2356 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U901  ( .A(
        \U1/keyexpantion/SB0/n2516 ), .B(\U1/keyexpantion/SB0/n2477 ), .Y(
        \U1/keyexpantion/SB0/n2304 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U900  ( .A(
        \U1/keyexpantion/SB0/n2506 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2380 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U899  ( .A(
        \U1/keyexpantion/SB0/n2234 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2205 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U898  ( .A(
        \U1/keyexpantion/SB0/n2356 ), .B(\U1/keyexpantion/SB0/n2304 ), .C(
        \U1/keyexpantion/SB0/n2380 ), .D(\U1/keyexpantion/SB0/n2205 ), .Y(
        \U1/keyexpantion/SB0/n2145 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U897  ( .A(\U1/keyexpantion/SB0/n2148 ), 
        .B(\U1/keyexpantion/SB0/n2147 ), .C(\U1/keyexpantion/SB0/n2146 ), .D(
        \U1/keyexpantion/SB0/n2145 ), .Y(\U1/keyexpantion/SB0/n2191 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U896  ( .A(\U1/keyexpantion/SB0/n2183 ), 
        .B(\U1/keyexpantion/SB0/n2202 ), .C(\U1/keyexpantion/SB0/n2529 ), .D(
        \U1/keyexpantion/SB0/n2191 ), .Y(\U1/keyexpantion/SB0/n2158 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U895  ( .A(\U1/keyexpantion/SB0/n2483 ), 
        .Y(\U1/keyexpantion/SB0/n2407 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U894  ( .A0(
        \U1/keyexpantion/SB0/n2359 ), .A1(\U1/keyexpantion/SB0/n2165 ), .B0(
        \U1/keyexpantion/SB0/n2303 ), .B1(\U1/keyexpantion/SB0/n2514 ), .Y(
        \U1/keyexpantion/SB0/n2149 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U893  ( .A0(
        \U1/keyexpantion/SB0/n2407 ), .A1(\U1/keyexpantion/SB0/n2459 ), .B0(
        \U1/keyexpantion/SB0/n2508 ), .B1(\U1/keyexpantion/SB0/n2516 ), .C0(
        \U1/keyexpantion/SB0/n2149 ), .Y(\U1/keyexpantion/SB0/n2157 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U892  ( .A(
        \U1/keyexpantion/SB0/n2428 ), .B(\U1/keyexpantion/SB0/n2431 ), .Y(
        \U1/keyexpantion/SB0/n2427 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U891  ( .A0(
        \U1/keyexpantion/SB0/n2362 ), .A1(\U1/keyexpantion/SB0/n2431 ), .B0(
        \U1/keyexpantion/SB0/n2319 ), .B1(\U1/keyexpantion/SB0/n2472 ), .Y(
        \U1/keyexpantion/SB0/n2150 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U890  ( .A0(
        \U1/keyexpantion/SB0/n2234 ), .A1(\U1/keyexpantion/SB0/n2427 ), .B0(
        \U1/keyexpantion/SB0/n2478 ), .B1(\U1/keyexpantion/SB0/n2497 ), .C0(
        \U1/keyexpantion/SB0/n2150 ), .Y(\U1/keyexpantion/SB0/n2156 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U889  ( .A(
        \U1/keyexpantion/SB0/n2502 ), .B(\U1/keyexpantion/SB0/n2361 ), .Y(
        \U1/keyexpantion/SB0/n2154 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U888  ( .A(\U1/keyexpantion/SB0/n2452 ), .B(\U1/keyexpantion/SB0/n2477 ), .Y(\U1/keyexpantion/SB0/n2419 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U887  ( .A(\U1/keyexpantion/SB0/n2419 ), 
        .Y(\U1/keyexpantion/SB0/n2153 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U886  ( .A(\U1/keyexpantion/SB0/n2410 ), .B(\U1/keyexpantion/SB0/n2483 ), .Y(\U1/keyexpantion/SB0/n2266 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U885  ( .A(\U1/keyexpantion/SB0/n2488 ), .B(\U1/keyexpantion/SB0/n2486 ), .Y(\U1/keyexpantion/SB0/n2444 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U884  ( .A(\U1/keyexpantion/SB0/n2444 ), 
        .Y(\U1/keyexpantion/SB0/n2151 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U883  ( .A(
        \U1/keyexpantion/SB0/n2459 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2276 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U882  ( .AN(
        \U1/keyexpantion/SB0/n2266 ), .B(\U1/keyexpantion/SB0/n2151 ), .C(
        \U1/keyexpantion/SB0/n2276 ), .Y(\U1/keyexpantion/SB0/n2152 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U881  ( .A0(
        \U1/keyexpantion/SB0/n2418 ), .A1(\U1/keyexpantion/SB0/n2154 ), .B0(
        \U1/keyexpantion/SB0/n2395 ), .B1(\U1/keyexpantion/SB0/n2153 ), .C0(
        \U1/keyexpantion/SB0/n2152 ), .Y(\U1/keyexpantion/SB0/n2155 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U880  ( .AN(
        \U1/keyexpantion/SB0/n2158 ), .B(\U1/keyexpantion/SB0/n2157 ), .C(
        \U1/keyexpantion/SB0/n2156 ), .D(\U1/keyexpantion/SB0/n2155 ), .Y(
        \U1/keyexpantion/ws [16]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U879  ( .A(\U1/keyexpantion/SB0/n2431 ), .B(\U1/keyexpantion/SB0/n2223 ), .Y(\U1/keyexpantion/SB0/n2283 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U878  ( .A(\U1/keyexpantion/SB0/n2378 ), .B(\U1/keyexpantion/SB0/n2428 ), .Y(\U1/keyexpantion/SB0/n2243 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U877  ( .A(\U1/keyexpantion/SB0/n2395 ), .B(\U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2377 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U876  ( .A0(
        \U1/keyexpantion/SB0/n2377 ), .A1(\U1/keyexpantion/SB0/n2431 ), .B0(
        \U1/keyexpantion/SB0/n2520 ), .Y(\U1/keyexpantion/SB0/n2163 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U875  ( .A(
        \U1/keyexpantion/SB0/n2459 ), .B(\U1/keyexpantion/SB0/n2507 ), .Y(
        \U1/keyexpantion/SB0/n2259 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U874  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2459 ), .Y(
        \U1/keyexpantion/SB0/n2383 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U873  ( .A(
        \U1/keyexpantion/SB0/n2504 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2291 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U872  ( .A(
        \U1/keyexpantion/SB0/n2259 ), .B(\U1/keyexpantion/SB0/n2383 ), .C(
        \U1/keyexpantion/SB0/n2291 ), .Y(\U1/keyexpantion/SB0/n2162 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U871  ( .A(\U1/keyexpantion/SB0/n2459 ), .B(\U1/keyexpantion/SB0/n2518 ), .Y(\U1/keyexpantion/SB0/n2318 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U870  ( .A(\U1/keyexpantion/SB0/n2504 ), .B(\U1/keyexpantion/SB0/n2495 ), .C(\U1/keyexpantion/SB0/n2516 ), .Y(
        \U1/keyexpantion/SB0/n2159 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U869  ( .A0(
        \U1/keyexpantion/SB0/n2318 ), .A1(\U1/keyexpantion/SB0/n2484 ), .B0(
        \U1/keyexpantion/SB0/n2159 ), .B1(\U1/keyexpantion/SB0/n2514 ), .C0(
        \U1/keyexpantion/SB0/n2378 ), .C1(\U1/keyexpantion/SB0/n2410 ), .Y(
        \U1/keyexpantion/SB0/n2161 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U868  ( .A0(
        \U1/keyexpantion/SB0/n2485 ), .A1(\U1/keyexpantion/SB0/n2513 ), .B0(
        \U1/keyexpantion/SB0/n2486 ), .B1(\U1/keyexpantion/SB0/n2483 ), .Y(
        \U1/keyexpantion/SB0/n2160 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U867  ( .A(\U1/keyexpantion/SB0/n2283 ), 
        .B(\U1/keyexpantion/SB0/n2243 ), .C(\U1/keyexpantion/SB0/n2163 ), .D(
        \U1/keyexpantion/SB0/n2162 ), .E(\U1/keyexpantion/SB0/n2161 ), .F(
        \U1/keyexpantion/SB0/n2160 ), .Y(\U1/keyexpantion/SB0/n2528 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U866  ( .A(\U1/keyexpantion/SB0/n2359 ), .B(\U1/keyexpantion/SB0/n2319 ), .Y(\U1/keyexpantion/SB0/n2209 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U865  ( .A0(
        \U1/keyexpantion/SB0/n2359 ), .A1(\U1/keyexpantion/SB0/n2449 ), .B0(
        \U1/keyexpantion/SB0/n2223 ), .Y(\U1/keyexpantion/SB0/n2170 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U864  ( .A(\U1/keyexpantion/SB0/n2453 ), .B(\U1/keyexpantion/SB0/n2459 ), .Y(\U1/keyexpantion/SB0/n2211 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U863  ( .A0(
        \U1/keyexpantion/SB0/n2316 ), .A1(\U1/keyexpantion/SB0/n2488 ), .B0(
        \U1/keyexpantion/SB0/n2211 ), .B1(\U1/keyexpantion/SB0/n2502 ), .Y(
        \U1/keyexpantion/SB0/n2169 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U862  ( .A0(
        \U1/keyexpantion/SB0/n2303 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2472 ), .B1(\U1/keyexpantion/SB0/n2378 ), .C0(
        \U1/keyexpantion/SB0/n2486 ), .C1(\U1/keyexpantion/SB0/n2429 ), .Y(
        \U1/keyexpantion/SB0/n2168 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U861  ( .A(\U1/keyexpantion/SB0/n2521 ), .B(\U1/keyexpantion/SB0/n2164 ), .Y(\U1/keyexpantion/SB0/n2267 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U860  ( .A(
        \U1/keyexpantion/SB0/n2508 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2274 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U859  ( .A(
        \U1/keyexpantion/SB0/n2450 ), .B(\U1/keyexpantion/SB0/n2503 ), .Y(
        \U1/keyexpantion/SB0/n2284 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U858  ( .A(
        \U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2518 ), .Y(
        \U1/keyexpantion/SB0/n2413 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U857  ( .AN(
        \U1/keyexpantion/SB0/n2267 ), .B(\U1/keyexpantion/SB0/n2274 ), .C(
        \U1/keyexpantion/SB0/n2284 ), .D(\U1/keyexpantion/SB0/n2413 ), .Y(
        \U1/keyexpantion/SB0/n2167 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U856  ( .A(\U1/keyexpantion/SB0/n2410 ), .B(\U1/keyexpantion/SB0/n2165 ), .Y(\U1/keyexpantion/SB0/n2392 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U855  ( .A(\U1/keyexpantion/SB0/n2488 ), .B(\U1/keyexpantion/SB0/n2472 ), .Y(\U1/keyexpantion/SB0/n2445 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U853  ( .A(
        \U1/keyexpantion/SB0/n2208 ), .B(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2233 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U851  ( .A(\U1/keyexpantion/SB0/n2209 ), 
        .B(\U1/keyexpantion/SB0/n2170 ), .C(\U1/keyexpantion/SB0/n2169 ), .D(
        \U1/keyexpantion/SB0/n2168 ), .E(\U1/keyexpantion/SB0/n2167 ), .F(
        \U1/keyexpantion/SB0/n2166 ), .Y(\U1/keyexpantion/SB0/n2203 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U850  ( .A(\U1/keyexpantion/SB0/n2426 ), .B(\U1/keyexpantion/SB0/n2223 ), .Y(\U1/keyexpantion/SB0/n2221 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U849  ( .A(\U1/keyexpantion/SB0/n2378 ), .B(\U1/keyexpantion/SB0/n2303 ), .Y(\U1/keyexpantion/SB0/n2458 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U848  ( .A(\U1/keyexpantion/SB0/n2359 ), .B(\U1/keyexpantion/SB0/n2429 ), .Y(\U1/keyexpantion/SB0/n2271 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U847  ( .A(\U1/keyexpantion/SB0/n2523 ), .B(\U1/keyexpantion/SB0/n2429 ), .Y(\U1/keyexpantion/SB0/n2286 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U846  ( .A(
        \U1/keyexpantion/SB0/n2454 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2371 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U845  ( .A(
        \U1/keyexpantion/SB0/n2504 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2238 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U844  ( .A(
        \U1/keyexpantion/SB0/n2508 ), .B(\U1/keyexpantion/SB0/n2504 ), .Y(
        \U1/keyexpantion/SB0/n2357 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U843  ( .A(
        \U1/keyexpantion/SB0/n2418 ), .B(\U1/keyexpantion/SB0/n2475 ), .Y(
        \U1/keyexpantion/SB0/n2257 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U842  ( .A(
        \U1/keyexpantion/SB0/n2371 ), .B(\U1/keyexpantion/SB0/n2238 ), .C(
        \U1/keyexpantion/SB0/n2357 ), .D(\U1/keyexpantion/SB0/n2257 ), .Y(
        \U1/keyexpantion/SB0/n2174 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U841  ( .A(\U1/keyexpantion/SB0/n2523 ), .B(\U1/keyexpantion/SB0/n2319 ), .Y(\U1/keyexpantion/SB0/n2307 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U840  ( .A(\U1/keyexpantion/SB0/n2522 ), .B(\U1/keyexpantion/SB0/n2303 ), .Y(\U1/keyexpantion/SB0/n2432 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U839  ( .A(\U1/keyexpantion/SB0/n2449 ), .B(\U1/keyexpantion/SB0/n2488 ), .Y(\U1/keyexpantion/SB0/n2382 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U838  ( .A(\U1/keyexpantion/SB0/n2410 ), .B(\U1/keyexpantion/SB0/n2488 ), .Y(\U1/keyexpantion/SB0/n2207 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U837  ( .A0(
        \U1/keyexpantion/SB0/n2488 ), .A1(\U1/keyexpantion/SB0/n2523 ), .B0(
        \U1/keyexpantion/SB0/n2319 ), .B1(\U1/keyexpantion/SB0/n2449 ), .Y(
        \U1/keyexpantion/SB0/n2172 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U836  ( .A0(
        \U1/keyexpantion/SB0/n2303 ), .A1(\U1/keyexpantion/SB0/n2520 ), .B0(
        \U1/keyexpantion/SB0/n2316 ), .B1(\U1/keyexpantion/SB0/n2378 ), .Y(
        \U1/keyexpantion/SB0/n2171 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U835  ( .A(\U1/keyexpantion/SB0/n2307 ), 
        .B(\U1/keyexpantion/SB0/n2432 ), .C(\U1/keyexpantion/SB0/n2382 ), .D(
        \U1/keyexpantion/SB0/n2207 ), .E(\U1/keyexpantion/SB0/n2172 ), .F(
        \U1/keyexpantion/SB0/n2171 ), .Y(\U1/keyexpantion/SB0/n2173 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U834  ( .A(\U1/keyexpantion/SB0/n2221 ), 
        .B(\U1/keyexpantion/SB0/n2458 ), .C(\U1/keyexpantion/SB0/n2271 ), .D(
        \U1/keyexpantion/SB0/n2286 ), .E(\U1/keyexpantion/SB0/n2174 ), .F(
        \U1/keyexpantion/SB0/n2173 ), .Y(\U1/keyexpantion/SB0/n2192 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U833  ( .A0(
        \U1/keyexpantion/SB0/n2454 ), .A1(\U1/keyexpantion/SB0/n2451 ), .B0(
        \U1/keyexpantion/SB0/n2507 ), .B1(\U1/keyexpantion/SB0/n2395 ), .C0(
        \U1/keyexpantion/SB0/n2192 ), .Y(\U1/keyexpantion/SB0/n2175 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U832  ( .A(\U1/keyexpantion/SB0/n2175 ), 
        .Y(\U1/keyexpantion/SB0/n2182 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U831  ( .A(
        \U1/keyexpantion/SB0/n2486 ), .B(\U1/keyexpantion/SB0/n2449 ), .Y(
        \U1/keyexpantion/SB0/n2476 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U830  ( .A0(
        \U1/keyexpantion/SB0/n2453 ), .A1(\U1/keyexpantion/SB0/n2476 ), .B0(
        \U1/keyexpantion/SB0/n2508 ), .Y(\U1/keyexpantion/SB0/n2178 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U829  ( .A0(
        \U1/keyexpantion/SB0/n2418 ), .A1(\U1/keyexpantion/SB0/n2497 ), .B0(
        \U1/keyexpantion/SB0/n2460 ), .Y(\U1/keyexpantion/SB0/n2177 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U828  ( .A0(
        \U1/keyexpantion/SB0/n2417 ), .A1(\U1/keyexpantion/SB0/n2459 ), .B0(
        \U1/keyexpantion/SB0/n2503 ), .Y(\U1/keyexpantion/SB0/n2176 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U827  ( .A(
        \U1/keyexpantion/SB0/n2450 ), .B(\U1/keyexpantion/SB0/n2496 ), .Y(
        \U1/keyexpantion/SB0/n2250 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U826  ( .A(
        \U1/keyexpantion/SB0/n2178 ), .B(\U1/keyexpantion/SB0/n2177 ), .C(
        \U1/keyexpantion/SB0/n2176 ), .D(\U1/keyexpantion/SB0/n2250 ), .Y(
        \U1/keyexpantion/SB0/n2181 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U825  ( .A(\U1/keyexpantion/SB0/n2495 ), .B(\U1/keyexpantion/SB0/n2411 ), .Y(\U1/keyexpantion/SB0/n2465 ) );
  AND3_X0P5M_A12TL \U1/keyexpantion/SB0/U824  ( .A(\U1/keyexpantion/SB0/n2465 ), .B(\U1/keyexpantion/SB0/n2485 ), .C(\U1/keyexpantion/SB0/n2472 ), .Y(
        \U1/keyexpantion/SB0/n2179 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U823  ( .A0(
        \U1/keyexpantion/SB0/n2449 ), .A1(\U1/keyexpantion/SB0/n2522 ), .B0(
        \U1/keyexpantion/SB0/n2179 ), .B1(\U1/keyexpantion/SB0/n2483 ), .C0(
        \U1/keyexpantion/SB0/n2521 ), .C1(\U1/keyexpantion/SB0/n2513 ), .Y(
        \U1/keyexpantion/SB0/n2180 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U822  ( .A(\U1/keyexpantion/SB0/n2528 ), 
        .B(\U1/keyexpantion/SB0/n2203 ), .C(\U1/keyexpantion/SB0/n2183 ), .D(
        \U1/keyexpantion/SB0/n2182 ), .E(\U1/keyexpantion/SB0/n2181 ), .F(
        \U1/keyexpantion/SB0/n2180 ), .Y(\U1/keyexpantion/ws [17]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U821  ( .A0(
        \U1/keyexpantion/SB0/n2477 ), .A1(\U1/keyexpantion/SB0/n2497 ), .B0(
        \U1/keyexpantion/SB0/n2518 ), .B1(\U1/keyexpantion/SB0/n2508 ), .Y(
        \U1/keyexpantion/SB0/n2184 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U820  ( .A0(
        \U1/keyexpantion/SB0/n2428 ), .A1(\U1/keyexpantion/SB0/n2522 ), .B0(
        \U1/keyexpantion/SB0/n2378 ), .B1(\U1/keyexpantion/SB0/n2449 ), .C0(
        \U1/keyexpantion/SB0/n2184 ), .Y(\U1/keyexpantion/SB0/n2190 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U819  ( .A(
        \U1/keyexpantion/SB0/n2503 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2287 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U818  ( .A(
        \U1/keyexpantion/SB0/n2477 ), .B(\U1/keyexpantion/SB0/n2453 ), .Y(
        \U1/keyexpantion/SB0/n2268 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U817  ( .A(
        \U1/keyexpantion/SB0/n2497 ), .B(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2236 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U816  ( .A(
        \U1/keyexpantion/SB0/n2417 ), .B(\U1/keyexpantion/SB0/n2460 ), .Y(
        \U1/keyexpantion/SB0/n2255 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U815  ( .A(
        \U1/keyexpantion/SB0/n2287 ), .B(\U1/keyexpantion/SB0/n2268 ), .C(
        \U1/keyexpantion/SB0/n2236 ), .D(\U1/keyexpantion/SB0/n2255 ), .Y(
        \U1/keyexpantion/SB0/n2189 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U814  ( .A(
        \U1/keyexpantion/SB0/n2523 ), .B(\U1/keyexpantion/SB0/n2501 ), .Y(
        \U1/keyexpantion/SB0/n2406 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U813  ( .A0(
        \U1/keyexpantion/SB0/n2454 ), .A1(\U1/keyexpantion/SB0/n2406 ), .B0(
        \U1/keyexpantion/SB0/n2507 ), .Y(\U1/keyexpantion/SB0/n2187 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U812  ( .A0(
        \U1/keyexpantion/SB0/n2504 ), .A1(\U1/keyexpantion/SB0/n2395 ), .B0(
        \U1/keyexpantion/SB0/n2407 ), .Y(\U1/keyexpantion/SB0/n2186 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U811  ( .A0(
        \U1/keyexpantion/SB0/n2412 ), .A1(\U1/keyexpantion/SB0/n2452 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2185 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U810  ( .A(
        \U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2504 ), .Y(
        \U1/keyexpantion/SB0/n2379 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U809  ( .A(
        \U1/keyexpantion/SB0/n2187 ), .B(\U1/keyexpantion/SB0/n2186 ), .C(
        \U1/keyexpantion/SB0/n2185 ), .D(\U1/keyexpantion/SB0/n2379 ), .Y(
        \U1/keyexpantion/SB0/n2188 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U808  ( .A(\U1/keyexpantion/SB0/n2193 ), 
        .B(\U1/keyexpantion/SB0/n2192 ), .C(\U1/keyexpantion/SB0/n2191 ), .D(
        \U1/keyexpantion/SB0/n2190 ), .E(\U1/keyexpantion/SB0/n2189 ), .F(
        \U1/keyexpantion/SB0/n2188 ), .Y(\U1/keyexpantion/SB0/n2527 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U807  ( .A0(
        \U1/keyexpantion/SB0/n2308 ), .A1(\U1/keyexpantion/SB0/n2508 ), .B0(
        \U1/keyexpantion/SB0/n2516 ), .B1(\U1/keyexpantion/SB0/n2451 ), .C0(
        \U1/keyexpantion/SB0/n2527 ), .Y(\U1/keyexpantion/SB0/n2194 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U806  ( .A(\U1/keyexpantion/SB0/n2194 ), 
        .Y(\U1/keyexpantion/SB0/n2201 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U805  ( .A(\U1/keyexpantion/SB0/n2460 ), .B(\U1/keyexpantion/SB0/n2222 ), .Y(\U1/keyexpantion/SB0/n2369 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U804  ( .A1N(
        \U1/keyexpantion/SB0/n2369 ), .A0(\U1/keyexpantion/SB0/n2478 ), .B0(
        \U1/keyexpantion/SB0/n2450 ), .Y(\U1/keyexpantion/SB0/n2197 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U803  ( .A0(
        \U1/keyexpantion/SB0/n2418 ), .A1(\U1/keyexpantion/SB0/n2301 ), .B0(
        \U1/keyexpantion/SB0/n2477 ), .Y(\U1/keyexpantion/SB0/n2196 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U802  ( .A0(
        \U1/keyexpantion/SB0/n2504 ), .A1(\U1/keyexpantion/SB0/n2459 ), .B0(
        \U1/keyexpantion/SB0/n2498 ), .Y(\U1/keyexpantion/SB0/n2195 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U801  ( .A(
        \U1/keyexpantion/SB0/n2475 ), .B(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2251 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U800  ( .A(
        \U1/keyexpantion/SB0/n2197 ), .B(\U1/keyexpantion/SB0/n2196 ), .C(
        \U1/keyexpantion/SB0/n2195 ), .D(\U1/keyexpantion/SB0/n2251 ), .Y(
        \U1/keyexpantion/SB0/n2200 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U799  ( .A(\U1/keyexpantion/SB0/n2474 ), .B(\U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2505 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U798  ( .A(\U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2452 ), .Y(\U1/keyexpantion/SB0/n2198 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U797  ( .A0(
        \U1/keyexpantion/SB0/n2505 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2198 ), .B1(\U1/keyexpantion/SB0/n2486 ), .C0(
        \U1/keyexpantion/SB0/n2429 ), .C1(\U1/keyexpantion/SB0/n2431 ), .Y(
        \U1/keyexpantion/SB0/n2199 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U796  ( .A(\U1/keyexpantion/SB0/n2204 ), 
        .B(\U1/keyexpantion/SB0/n2203 ), .C(\U1/keyexpantion/SB0/n2202 ), .D(
        \U1/keyexpantion/SB0/n2201 ), .E(\U1/keyexpantion/SB0/n2200 ), .F(
        \U1/keyexpantion/SB0/n2199 ), .Y(\U1/keyexpantion/ws [18]) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U795  ( .A(
        \U1/keyexpantion/SB0/n2308 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2510 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U794  ( .AN(
        \U1/keyexpantion/SB0/n2207 ), .B(\U1/keyexpantion/SB0/n2206 ), .C(
        \U1/keyexpantion/SB0/n2205 ), .D(\U1/keyexpantion/SB0/n2510 ), .Y(
        \U1/keyexpantion/SB0/n2214 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U793  ( .A0(
        \U1/keyexpantion/SB0/n2208 ), .A1(\U1/keyexpantion/SB0/n2477 ), .B0(
        \U1/keyexpantion/SB0/n2395 ), .Y(\U1/keyexpantion/SB0/n2210 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U790  ( .A(\U1/keyexpantion/SB0/n2451 ), .B(\U1/keyexpantion/SB0/n2498 ), .Y(\U1/keyexpantion/SB0/n2462 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U789  ( .A0(
        \U1/keyexpantion/SB0/n2316 ), .A1(\U1/keyexpantion/SB0/n2520 ), .B0(
        \U1/keyexpantion/SB0/n2462 ), .B1(\U1/keyexpantion/SB0/n2473 ), .C0(
        \U1/keyexpantion/SB0/n2514 ), .C1(\U1/keyexpantion/SB0/n2523 ), .Y(
        \U1/keyexpantion/SB0/n2212 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U788  ( .A(\U1/keyexpantion/SB0/n2217 ), 
        .B(\U1/keyexpantion/SB0/n2216 ), .C(\U1/keyexpantion/SB0/n2215 ), .D(
        \U1/keyexpantion/SB0/n2214 ), .E(\U1/keyexpantion/SB0/n2213 ), .F(
        \U1/keyexpantion/SB0/n2212 ), .Y(\U1/keyexpantion/SB0/n2425 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U787  ( .AN(
        \U1/keyexpantion/SB0/n2221 ), .B(\U1/keyexpantion/SB0/n2220 ), .C(
        \U1/keyexpantion/SB0/n2219 ), .D(\U1/keyexpantion/SB0/n2218 ), .Y(
        \U1/keyexpantion/SB0/n2231 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U786  ( .A0(
        \U1/keyexpantion/SB0/n2508 ), .A1(\U1/keyexpantion/SB0/n2418 ), .B0(
        \U1/keyexpantion/SB0/n2503 ), .B1(\U1/keyexpantion/SB0/n2417 ), .C0(
        \U1/keyexpantion/SB0/n2222 ), .C1(\U1/keyexpantion/SB0/n2518 ), .Y(
        \U1/keyexpantion/SB0/n2230 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U785  ( .A0(
        \U1/keyexpantion/SB0/n2472 ), .A1(\U1/keyexpantion/SB0/n2378 ), .B0(
        \U1/keyexpantion/SB0/n2223 ), .B1(\U1/keyexpantion/SB0/n2316 ), .Y(
        \U1/keyexpantion/SB0/n2224 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U784  ( .A0(
        \U1/keyexpantion/SB0/n2395 ), .A1(\U1/keyexpantion/SB0/n2412 ), .B0(
        \U1/keyexpantion/SB0/n2411 ), .B1(\U1/keyexpantion/SB0/n2475 ), .C0(
        \U1/keyexpantion/SB0/n2224 ), .Y(\U1/keyexpantion/SB0/n2229 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U783  ( .A(
        \U1/keyexpantion/SB0/n2483 ), .B(\U1/keyexpantion/SB0/n2522 ), .Y(
        \U1/keyexpantion/SB0/n2226 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U782  ( .A0(
        \U1/keyexpantion/SB0/n2308 ), .A1(\U1/keyexpantion/SB0/n2227 ), .B0(
        \U1/keyexpantion/SB0/n2504 ), .B1(\U1/keyexpantion/SB0/n2226 ), .C0(
        \U1/keyexpantion/SB0/n2225 ), .Y(\U1/keyexpantion/SB0/n2228 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U781  ( .AN(
        \U1/keyexpantion/SB0/n2231 ), .B(\U1/keyexpantion/SB0/n2230 ), .C(
        \U1/keyexpantion/SB0/n2229 ), .D(\U1/keyexpantion/SB0/n2228 ), .Y(
        \U1/keyexpantion/SB0/n2470 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U780  ( .A(\U1/keyexpantion/SB0/n2232 ), 
        .Y(\U1/keyexpantion/SB0/n2248 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U779  ( .A0(
        \U1/keyexpantion/SB0/n2362 ), .A1(\U1/keyexpantion/SB0/n2431 ), .B0(
        \U1/keyexpantion/SB0/n2233 ), .Y(\U1/keyexpantion/SB0/n2247 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U778  ( .A0(
        \U1/keyexpantion/SB0/n2504 ), .A1(\U1/keyexpantion/SB0/n2503 ), .B0(
        \U1/keyexpantion/SB0/n2474 ), .B1(\U1/keyexpantion/SB0/n2234 ), .Y(
        \U1/keyexpantion/SB0/n2235 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U777  ( .A0(
        \U1/keyexpantion/SB0/n2485 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2501 ), .B1(\U1/keyexpantion/SB0/n2513 ), .C0(
        \U1/keyexpantion/SB0/n2235 ), .Y(\U1/keyexpantion/SB0/n2246 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U776  ( .A(
        \U1/keyexpantion/SB0/n2239 ), .B(\U1/keyexpantion/SB0/n2238 ), .C(
        \U1/keyexpantion/SB0/n2237 ), .D(\U1/keyexpantion/SB0/n2236 ), .Y(
        \U1/keyexpantion/SB0/n2245 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U775  ( .AN(
        \U1/keyexpantion/SB0/n2243 ), .B(\U1/keyexpantion/SB0/n2242 ), .C(
        \U1/keyexpantion/SB0/n2241 ), .D(\U1/keyexpantion/SB0/n2240 ), .Y(
        \U1/keyexpantion/SB0/n2244 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U774  ( .A(\U1/keyexpantion/SB0/n2249 ), 
        .B(\U1/keyexpantion/SB0/n2248 ), .C(\U1/keyexpantion/SB0/n2247 ), .D(
        \U1/keyexpantion/SB0/n2246 ), .E(\U1/keyexpantion/SB0/n2245 ), .F(
        \U1/keyexpantion/SB0/n2244 ), .Y(\U1/keyexpantion/SB0/n2374 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U773  ( .A0(
        \U1/keyexpantion/SB0/n2461 ), .A1(\U1/keyexpantion/SB0/n2378 ), .B0(
        \U1/keyexpantion/SB0/n2250 ), .Y(\U1/keyexpantion/SB0/n2265 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U772  ( .AN(
        \U1/keyexpantion/SB0/n2254 ), .B(\U1/keyexpantion/SB0/n2253 ), .C(
        \U1/keyexpantion/SB0/n2252 ), .D(\U1/keyexpantion/SB0/n2251 ), .Y(
        \U1/keyexpantion/SB0/n2264 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U771  ( .A(
        \U1/keyexpantion/SB0/n2495 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2509 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U770  ( .A(
        \U1/keyexpantion/SB0/n2257 ), .B(\U1/keyexpantion/SB0/n2256 ), .C(
        \U1/keyexpantion/SB0/n2255 ), .D(\U1/keyexpantion/SB0/n2509 ), .Y(
        \U1/keyexpantion/SB0/n2263 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U769  ( .A(
        \U1/keyexpantion/SB0/n2261 ), .B(\U1/keyexpantion/SB0/n2260 ), .C(
        \U1/keyexpantion/SB0/n2259 ), .D(\U1/keyexpantion/SB0/n2258 ), .Y(
        \U1/keyexpantion/SB0/n2262 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U768  ( .A(\U1/keyexpantion/SB0/n2267 ), 
        .B(\U1/keyexpantion/SB0/n2266 ), .C(\U1/keyexpantion/SB0/n2265 ), .D(
        \U1/keyexpantion/SB0/n2264 ), .E(\U1/keyexpantion/SB0/n2263 ), .F(
        \U1/keyexpantion/SB0/n2262 ), .Y(\U1/keyexpantion/SB0/n2398 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U767  ( .AN(
        \U1/keyexpantion/SB0/n2271 ), .B(\U1/keyexpantion/SB0/n2270 ), .C(
        \U1/keyexpantion/SB0/n2269 ), .D(\U1/keyexpantion/SB0/n2268 ), .Y(
        \U1/keyexpantion/SB0/n2280 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U766  ( .A(
        \U1/keyexpantion/SB0/n2275 ), .B(\U1/keyexpantion/SB0/n2274 ), .C(
        \U1/keyexpantion/SB0/n2273 ), .D(\U1/keyexpantion/SB0/n2272 ), .Y(
        \U1/keyexpantion/SB0/n2279 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U765  ( .A(\U1/keyexpantion/SB0/n2460 ), .B(\U1/keyexpantion/SB0/n2496 ), .C(\U1/keyexpantion/SB0/n2498 ), .Y(
        \U1/keyexpantion/SB0/n2277 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U764  ( .A0(
        \U1/keyexpantion/SB0/n2277 ), .A1(\U1/keyexpantion/SB0/n2486 ), .B0(
        \U1/keyexpantion/SB0/n2316 ), .B1(\U1/keyexpantion/SB0/n2522 ), .C0(
        \U1/keyexpantion/SB0/n2276 ), .Y(\U1/keyexpantion/SB0/n2278 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U763  ( .A(\U1/keyexpantion/SB0/n2283 ), 
        .B(\U1/keyexpantion/SB0/n2282 ), .C(\U1/keyexpantion/SB0/n2281 ), .D(
        \U1/keyexpantion/SB0/n2280 ), .E(\U1/keyexpantion/SB0/n2279 ), .F(
        \U1/keyexpantion/SB0/n2278 ), .Y(\U1/keyexpantion/SB0/n2446 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U762  ( .A0(
        \U1/keyexpantion/SB0/n2316 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2284 ), .Y(\U1/keyexpantion/SB0/n2298 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U761  ( .A0(
        \U1/keyexpantion/SB0/n2450 ), .A1(\U1/keyexpantion/SB0/n2452 ), .B0(
        \U1/keyexpantion/SB0/n2507 ), .B1(\U1/keyexpantion/SB0/n2417 ), .Y(
        \U1/keyexpantion/SB0/n2285 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U760  ( .A0(
        \U1/keyexpantion/SB0/n2361 ), .A1(\U1/keyexpantion/SB0/n2449 ), .B0(
        \U1/keyexpantion/SB0/n2362 ), .B1(\U1/keyexpantion/SB0/n2426 ), .C0(
        \U1/keyexpantion/SB0/n2285 ), .Y(\U1/keyexpantion/SB0/n2297 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U759  ( .A(\U1/keyexpantion/SB0/n2286 ), 
        .Y(\U1/keyexpantion/SB0/n2289 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U758  ( .AN(
        \U1/keyexpantion/SB0/n2290 ), .B(\U1/keyexpantion/SB0/n2289 ), .C(
        \U1/keyexpantion/SB0/n2288 ), .D(\U1/keyexpantion/SB0/n2287 ), .Y(
        \U1/keyexpantion/SB0/n2296 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U757  ( .A(
        \U1/keyexpantion/SB0/n2294 ), .B(\U1/keyexpantion/SB0/n2293 ), .C(
        \U1/keyexpantion/SB0/n2292 ), .D(\U1/keyexpantion/SB0/n2291 ), .Y(
        \U1/keyexpantion/SB0/n2295 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U756  ( .A(\U1/keyexpantion/SB0/n2300 ), 
        .B(\U1/keyexpantion/SB0/n2299 ), .C(\U1/keyexpantion/SB0/n2298 ), .D(
        \U1/keyexpantion/SB0/n2297 ), .E(\U1/keyexpantion/SB0/n2296 ), .F(
        \U1/keyexpantion/SB0/n2295 ), .Y(\U1/keyexpantion/SB0/n2405 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U755  ( .A0(
        \U1/keyexpantion/SB0/n2496 ), .A1(\U1/keyexpantion/SB0/n2301 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .B1(\U1/keyexpantion/SB0/n2452 ), .Y(
        \U1/keyexpantion/SB0/n2302 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U754  ( .A0(
        \U1/keyexpantion/SB0/n2378 ), .A1(\U1/keyexpantion/SB0/n2523 ), .B0(
        \U1/keyexpantion/SB0/n2303 ), .B1(\U1/keyexpantion/SB0/n2513 ), .C0(
        \U1/keyexpantion/SB0/n2302 ), .Y(\U1/keyexpantion/SB0/n2315 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U753  ( .AN(
        \U1/keyexpantion/SB0/n2307 ), .B(\U1/keyexpantion/SB0/n2306 ), .C(
        \U1/keyexpantion/SB0/n2305 ), .D(\U1/keyexpantion/SB0/n2304 ), .Y(
        \U1/keyexpantion/SB0/n2314 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U752  ( .A0(
        \U1/keyexpantion/SB0/n2516 ), .A1(\U1/keyexpantion/SB0/n2308 ), .B0(
        \U1/keyexpantion/SB0/n2507 ), .Y(\U1/keyexpantion/SB0/n2312 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U751  ( .A(
        \U1/keyexpantion/SB0/n2483 ), .B(\U1/keyexpantion/SB0/n2488 ), .Y(
        \U1/keyexpantion/SB0/n2309 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U750  ( .A0(
        \U1/keyexpantion/SB0/n2459 ), .A1(\U1/keyexpantion/SB0/n2309 ), .B0(
        \U1/keyexpantion/SB0/n2460 ), .B1(\U1/keyexpantion/SB0/n2406 ), .Y(
        \U1/keyexpantion/SB0/n2310 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U749  ( .A(
        \U1/keyexpantion/SB0/n2312 ), .B(\U1/keyexpantion/SB0/n2311 ), .C(
        \U1/keyexpantion/SB0/n2310 ), .Y(\U1/keyexpantion/SB0/n2313 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U748  ( .A(\U1/keyexpantion/SB0/n2398 ), 
        .B(\U1/keyexpantion/SB0/n2446 ), .C(\U1/keyexpantion/SB0/n2405 ), .D(
        \U1/keyexpantion/SB0/n2315 ), .E(\U1/keyexpantion/SB0/n2314 ), .F(
        \U1/keyexpantion/SB0/n2313 ), .Y(\U1/keyexpantion/SB0/n2492 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U747  ( .A(\U1/keyexpantion/SB0/n2425 ), 
        .B(\U1/keyexpantion/SB0/n2470 ), .C(\U1/keyexpantion/SB0/n2374 ), .D(
        \U1/keyexpantion/SB0/n2492 ), .Y(\U1/keyexpantion/SB0/n2329 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U746  ( .A0(
        \U1/keyexpantion/SB0/n2472 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2316 ), .B1(\U1/keyexpantion/SB0/n2488 ), .Y(
        \U1/keyexpantion/SB0/n2317 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U745  ( .A0(
        \U1/keyexpantion/SB0/n2477 ), .A1(\U1/keyexpantion/SB0/n2495 ), .B0(
        \U1/keyexpantion/SB0/n2508 ), .B1(\U1/keyexpantion/SB0/n2516 ), .C0(
        \U1/keyexpantion/SB0/n2317 ), .Y(\U1/keyexpantion/SB0/n2328 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U744  ( .A(\U1/keyexpantion/SB0/n2318 ), 
        .Y(\U1/keyexpantion/SB0/n2321 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U743  ( .A0(
        \U1/keyexpantion/SB0/n2319 ), .A1(\U1/keyexpantion/SB0/n2449 ), .B0(
        \U1/keyexpantion/SB0/n2377 ), .B1(\U1/keyexpantion/SB0/n2429 ), .Y(
        \U1/keyexpantion/SB0/n2320 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U742  ( .A0(
        \U1/keyexpantion/SB0/n2496 ), .A1(\U1/keyexpantion/SB0/n2321 ), .B0(
        \U1/keyexpantion/SB0/n2478 ), .B1(\U1/keyexpantion/SB0/n2427 ), .C0(
        \U1/keyexpantion/SB0/n2320 ), .Y(\U1/keyexpantion/SB0/n2327 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U741  ( .A0(
        \U1/keyexpantion/SB0/n2518 ), .A1(\U1/keyexpantion/SB0/n2395 ), .B0(
        \U1/keyexpantion/SB0/n2498 ), .Y(\U1/keyexpantion/SB0/n2325 ) );
  AND4_X0P5M_A12TL \U1/keyexpantion/SB0/U740  ( .A(\U1/keyexpantion/SB0/n2325 ), .B(\U1/keyexpantion/SB0/n2324 ), .C(\U1/keyexpantion/SB0/n2323 ), .D(
        \U1/keyexpantion/SB0/n2322 ), .Y(\U1/keyexpantion/SB0/n2326 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U739  ( .AN(
        \U1/keyexpantion/SB0/n2329 ), .B(\U1/keyexpantion/SB0/n2328 ), .C(
        \U1/keyexpantion/SB0/n2327 ), .D(\U1/keyexpantion/SB0/n2326 ), .Y(
        \U1/keyexpantion/ws [19]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U738  ( .A(\U1/keyexpantion/SB0/n3175 ), .B(\U1/keyexpantion/SB0/n2992 ), .Y(\U1/keyexpantion/SB0/n3052 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U737  ( .A(\U1/keyexpantion/SB0/n3122 ), .B(\U1/keyexpantion/SB0/n3172 ), .Y(\U1/keyexpantion/SB0/n3012 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U736  ( .A(\U1/keyexpantion/SB0/n3139 ), .B(\U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n3121 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U735  ( .A0(
        \U1/keyexpantion/SB0/n3121 ), .A1(\U1/keyexpantion/SB0/n3175 ), .B0(
        \U1/keyexpantion/SB0/n3264 ), .Y(\U1/keyexpantion/SB0/n2334 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U734  ( .A(
        \U1/keyexpantion/SB0/n3203 ), .B(\U1/keyexpantion/SB0/n3251 ), .Y(
        \U1/keyexpantion/SB0/n3028 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U733  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3203 ), .Y(
        \U1/keyexpantion/SB0/n3127 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U732  ( .A(
        \U1/keyexpantion/SB0/n3248 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3060 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U731  ( .A(
        \U1/keyexpantion/SB0/n3028 ), .B(\U1/keyexpantion/SB0/n3127 ), .C(
        \U1/keyexpantion/SB0/n3060 ), .Y(\U1/keyexpantion/SB0/n2333 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U730  ( .A(\U1/keyexpantion/SB0/n3203 ), .B(\U1/keyexpantion/SB0/n3262 ), .Y(\U1/keyexpantion/SB0/n3087 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U729  ( .A(\U1/keyexpantion/SB0/n3248 ), .B(\U1/keyexpantion/SB0/n3239 ), .C(\U1/keyexpantion/SB0/n3260 ), .Y(
        \U1/keyexpantion/SB0/n2330 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U728  ( .A0(
        \U1/keyexpantion/SB0/n3087 ), .A1(\U1/keyexpantion/SB0/n3228 ), .B0(
        \U1/keyexpantion/SB0/n2330 ), .B1(\U1/keyexpantion/SB0/n3258 ), .C0(
        \U1/keyexpantion/SB0/n3122 ), .C1(\U1/keyexpantion/SB0/n3154 ), .Y(
        \U1/keyexpantion/SB0/n2332 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U727  ( .A0(
        \U1/keyexpantion/SB0/n3229 ), .A1(\U1/keyexpantion/SB0/n3257 ), .B0(
        \U1/keyexpantion/SB0/n3230 ), .B1(\U1/keyexpantion/SB0/n3227 ), .Y(
        \U1/keyexpantion/SB0/n2331 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U726  ( .A(\U1/keyexpantion/SB0/n3052 ), 
        .B(\U1/keyexpantion/SB0/n3012 ), .C(\U1/keyexpantion/SB0/n2334 ), .D(
        \U1/keyexpantion/SB0/n2333 ), .E(\U1/keyexpantion/SB0/n2332 ), .F(
        \U1/keyexpantion/SB0/n2331 ), .Y(\U1/keyexpantion/SB0/n3272 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U725  ( .A(\U1/keyexpantion/SB0/n3103 ), .B(\U1/keyexpantion/SB0/n3088 ), .Y(\U1/keyexpantion/SB0/n2978 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U724  ( .A0(
        \U1/keyexpantion/SB0/n3103 ), .A1(\U1/keyexpantion/SB0/n3193 ), .B0(
        \U1/keyexpantion/SB0/n2992 ), .Y(\U1/keyexpantion/SB0/n2341 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U723  ( .A(\U1/keyexpantion/SB0/n3197 ), .B(\U1/keyexpantion/SB0/n3203 ), .Y(\U1/keyexpantion/SB0/n2980 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U722  ( .A0(
        \U1/keyexpantion/SB0/n3085 ), .A1(\U1/keyexpantion/SB0/n3232 ), .B0(
        \U1/keyexpantion/SB0/n2980 ), .B1(\U1/keyexpantion/SB0/n3246 ), .Y(
        \U1/keyexpantion/SB0/n2340 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U721  ( .A0(
        \U1/keyexpantion/SB0/n3072 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n3216 ), .B1(\U1/keyexpantion/SB0/n3122 ), .C0(
        \U1/keyexpantion/SB0/n3230 ), .C1(\U1/keyexpantion/SB0/n3173 ), .Y(
        \U1/keyexpantion/SB0/n2339 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U720  ( .A(\U1/keyexpantion/SB0/n3265 ), .B(\U1/keyexpantion/SB0/n2335 ), .Y(\U1/keyexpantion/SB0/n3036 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U719  ( .A(
        \U1/keyexpantion/SB0/n3252 ), .B(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3043 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U718  ( .A(
        \U1/keyexpantion/SB0/n3194 ), .B(\U1/keyexpantion/SB0/n3247 ), .Y(
        \U1/keyexpantion/SB0/n3053 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U717  ( .A(
        \U1/keyexpantion/SB0/n3222 ), .B(\U1/keyexpantion/SB0/n3262 ), .Y(
        \U1/keyexpantion/SB0/n3157 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U716  ( .AN(
        \U1/keyexpantion/SB0/n3036 ), .B(\U1/keyexpantion/SB0/n3043 ), .C(
        \U1/keyexpantion/SB0/n3053 ), .D(\U1/keyexpantion/SB0/n3157 ), .Y(
        \U1/keyexpantion/SB0/n2338 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U715  ( .A(\U1/keyexpantion/SB0/n3154 ), .B(\U1/keyexpantion/SB0/n2336 ), .Y(\U1/keyexpantion/SB0/n3136 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U714  ( .A(\U1/keyexpantion/SB0/n3232 ), .B(\U1/keyexpantion/SB0/n3216 ), .Y(\U1/keyexpantion/SB0/n3189 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U712  ( .A(
        \U1/keyexpantion/SB0/n2977 ), .B(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3002 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U710  ( .A(\U1/keyexpantion/SB0/n2978 ), 
        .B(\U1/keyexpantion/SB0/n2341 ), .C(\U1/keyexpantion/SB0/n2340 ), .D(
        \U1/keyexpantion/SB0/n2339 ), .E(\U1/keyexpantion/SB0/n2338 ), .F(
        \U1/keyexpantion/SB0/n2337 ), .Y(\U1/keyexpantion/SB0/n2913 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U709  ( .A(\U1/keyexpantion/SB0/n3170 ), .B(\U1/keyexpantion/SB0/n2992 ), .Y(\U1/keyexpantion/SB0/n2990 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U708  ( .A(\U1/keyexpantion/SB0/n3122 ), .B(\U1/keyexpantion/SB0/n3072 ), .Y(\U1/keyexpantion/SB0/n3202 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U707  ( .A(\U1/keyexpantion/SB0/n3103 ), .B(\U1/keyexpantion/SB0/n3173 ), .Y(\U1/keyexpantion/SB0/n3040 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U706  ( .A(\U1/keyexpantion/SB0/n3267 ), .B(\U1/keyexpantion/SB0/n3173 ), .Y(\U1/keyexpantion/SB0/n3055 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U705  ( .A(
        \U1/keyexpantion/SB0/n3198 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3115 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U704  ( .A(
        \U1/keyexpantion/SB0/n3248 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3007 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U703  ( .A(
        \U1/keyexpantion/SB0/n3252 ), .B(\U1/keyexpantion/SB0/n3248 ), .Y(
        \U1/keyexpantion/SB0/n3101 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U702  ( .A(
        \U1/keyexpantion/SB0/n3162 ), .B(\U1/keyexpantion/SB0/n3219 ), .Y(
        \U1/keyexpantion/SB0/n3026 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U701  ( .A(
        \U1/keyexpantion/SB0/n3115 ), .B(\U1/keyexpantion/SB0/n3007 ), .C(
        \U1/keyexpantion/SB0/n3101 ), .D(\U1/keyexpantion/SB0/n3026 ), .Y(
        \U1/keyexpantion/SB0/n2345 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U700  ( .A(\U1/keyexpantion/SB0/n3267 ), .B(\U1/keyexpantion/SB0/n3088 ), .Y(\U1/keyexpantion/SB0/n3076 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U699  ( .A(\U1/keyexpantion/SB0/n3266 ), .B(\U1/keyexpantion/SB0/n3072 ), .Y(\U1/keyexpantion/SB0/n3176 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U698  ( .A(\U1/keyexpantion/SB0/n3193 ), .B(\U1/keyexpantion/SB0/n3232 ), .Y(\U1/keyexpantion/SB0/n3126 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U697  ( .A(\U1/keyexpantion/SB0/n3154 ), .B(\U1/keyexpantion/SB0/n3232 ), .Y(\U1/keyexpantion/SB0/n2976 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U696  ( .A0(
        \U1/keyexpantion/SB0/n3232 ), .A1(\U1/keyexpantion/SB0/n3267 ), .B0(
        \U1/keyexpantion/SB0/n3088 ), .B1(\U1/keyexpantion/SB0/n3193 ), .Y(
        \U1/keyexpantion/SB0/n2343 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U695  ( .A0(
        \U1/keyexpantion/SB0/n3072 ), .A1(\U1/keyexpantion/SB0/n3264 ), .B0(
        \U1/keyexpantion/SB0/n3085 ), .B1(\U1/keyexpantion/SB0/n3122 ), .Y(
        \U1/keyexpantion/SB0/n2342 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U694  ( .A(\U1/keyexpantion/SB0/n3076 ), 
        .B(\U1/keyexpantion/SB0/n3176 ), .C(\U1/keyexpantion/SB0/n3126 ), .D(
        \U1/keyexpantion/SB0/n2976 ), .E(\U1/keyexpantion/SB0/n2343 ), .F(
        \U1/keyexpantion/SB0/n2342 ), .Y(\U1/keyexpantion/SB0/n2344 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U693  ( .A(\U1/keyexpantion/SB0/n2990 ), 
        .B(\U1/keyexpantion/SB0/n3202 ), .C(\U1/keyexpantion/SB0/n3040 ), .D(
        \U1/keyexpantion/SB0/n3055 ), .E(\U1/keyexpantion/SB0/n2345 ), .F(
        \U1/keyexpantion/SB0/n2344 ), .Y(\U1/keyexpantion/SB0/n2902 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U692  ( .A0(
        \U1/keyexpantion/SB0/n3198 ), .A1(\U1/keyexpantion/SB0/n3195 ), .B0(
        \U1/keyexpantion/SB0/n3251 ), .B1(\U1/keyexpantion/SB0/n3139 ), .C0(
        \U1/keyexpantion/SB0/n2902 ), .Y(\U1/keyexpantion/SB0/n2346 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U691  ( .A(\U1/keyexpantion/SB0/n2346 ), 
        .Y(\U1/keyexpantion/SB0/n2353 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U690  ( .A(
        \U1/keyexpantion/SB0/n3230 ), .B(\U1/keyexpantion/SB0/n3193 ), .Y(
        \U1/keyexpantion/SB0/n3220 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U689  ( .A0(
        \U1/keyexpantion/SB0/n3197 ), .A1(\U1/keyexpantion/SB0/n3220 ), .B0(
        \U1/keyexpantion/SB0/n3252 ), .Y(\U1/keyexpantion/SB0/n2349 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U688  ( .A0(
        \U1/keyexpantion/SB0/n3162 ), .A1(\U1/keyexpantion/SB0/n3241 ), .B0(
        \U1/keyexpantion/SB0/n3204 ), .Y(\U1/keyexpantion/SB0/n2348 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U687  ( .A0(
        \U1/keyexpantion/SB0/n3161 ), .A1(\U1/keyexpantion/SB0/n3203 ), .B0(
        \U1/keyexpantion/SB0/n3247 ), .Y(\U1/keyexpantion/SB0/n2347 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U686  ( .A(
        \U1/keyexpantion/SB0/n3194 ), .B(\U1/keyexpantion/SB0/n3240 ), .Y(
        \U1/keyexpantion/SB0/n3019 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U685  ( .A(
        \U1/keyexpantion/SB0/n2349 ), .B(\U1/keyexpantion/SB0/n2348 ), .C(
        \U1/keyexpantion/SB0/n2347 ), .D(\U1/keyexpantion/SB0/n3019 ), .Y(
        \U1/keyexpantion/SB0/n2352 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U684  ( .A(\U1/keyexpantion/SB0/n3239 ), .B(\U1/keyexpantion/SB0/n3155 ), .Y(\U1/keyexpantion/SB0/n3209 ) );
  AND3_X0P5M_A12TL \U1/keyexpantion/SB0/U683  ( .A(\U1/keyexpantion/SB0/n3209 ), .B(\U1/keyexpantion/SB0/n3229 ), .C(\U1/keyexpantion/SB0/n3216 ), .Y(
        \U1/keyexpantion/SB0/n2350 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U682  ( .A0(
        \U1/keyexpantion/SB0/n3193 ), .A1(\U1/keyexpantion/SB0/n3266 ), .B0(
        \U1/keyexpantion/SB0/n2350 ), .B1(\U1/keyexpantion/SB0/n3227 ), .C0(
        \U1/keyexpantion/SB0/n3265 ), .C1(\U1/keyexpantion/SB0/n3257 ), .Y(
        \U1/keyexpantion/SB0/n2351 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U681  ( .A(\U1/keyexpantion/SB0/n3272 ), 
        .B(\U1/keyexpantion/SB0/n2913 ), .C(\U1/keyexpantion/SB0/n2354 ), .D(
        \U1/keyexpantion/SB0/n2353 ), .E(\U1/keyexpantion/SB0/n2352 ), .F(
        \U1/keyexpantion/SB0/n2351 ), .Y(\U1/keyexpantion/ws [1]) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U680  ( .A0(
        \U1/keyexpantion/SB0/n2369 ), .A1(\U1/keyexpantion/SB0/n2484 ), .B0(
        \U1/keyexpantion/SB0/n2428 ), .Y(\U1/keyexpantion/SB0/n2366 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U679  ( .A(
        \U1/keyexpantion/SB0/n2357 ), .B(\U1/keyexpantion/SB0/n2356 ), .C(
        \U1/keyexpantion/SB0/n2355 ), .Y(\U1/keyexpantion/SB0/n2365 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U678  ( .A(\U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2507 ), .Y(\U1/keyexpantion/SB0/n2360 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U677  ( .A(\U1/keyexpantion/SB0/n2478 ), .B(\U1/keyexpantion/SB0/n2412 ), .Y(\U1/keyexpantion/SB0/n2358 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U676  ( .A0(
        \U1/keyexpantion/SB0/n2360 ), .A1(\U1/keyexpantion/SB0/n2359 ), .B0(
        \U1/keyexpantion/SB0/n2358 ), .B1(\U1/keyexpantion/SB0/n2501 ), .C0(
        \U1/keyexpantion/SB0/n2484 ), .C1(\U1/keyexpantion/SB0/n2410 ), .Y(
        \U1/keyexpantion/SB0/n2364 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U675  ( .A0(
        \U1/keyexpantion/SB0/n2461 ), .A1(\U1/keyexpantion/SB0/n2362 ), .B0(
        \U1/keyexpantion/SB0/n2523 ), .B1(\U1/keyexpantion/SB0/n2513 ), .C0(
        \U1/keyexpantion/SB0/n2486 ), .C1(\U1/keyexpantion/SB0/n2361 ), .Y(
        \U1/keyexpantion/SB0/n2363 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U674  ( .A(\U1/keyexpantion/SB0/n2368 ), 
        .B(\U1/keyexpantion/SB0/n2367 ), .C(\U1/keyexpantion/SB0/n2366 ), .D(
        \U1/keyexpantion/SB0/n2365 ), .E(\U1/keyexpantion/SB0/n2364 ), .F(
        \U1/keyexpantion/SB0/n2363 ), .Y(\U1/keyexpantion/SB0/n2493 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U673  ( .A0(
        \U1/keyexpantion/SB0/n2369 ), .A1(\U1/keyexpantion/SB0/n2378 ), .B0(
        \U1/keyexpantion/SB0/n2449 ), .Y(\U1/keyexpantion/SB0/n2404 ) );
  AOI31_X0P5M_A12TL \U1/keyexpantion/SB0/U672  ( .A0(
        \U1/keyexpantion/SB0/n2473 ), .A1(\U1/keyexpantion/SB0/n2486 ), .A2(
        \U1/keyexpantion/SB0/n2426 ), .B0(\U1/keyexpantion/SB0/n2502 ), .Y(
        \U1/keyexpantion/SB0/n2403 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U671  ( .A(
        \U1/keyexpantion/SB0/n2373 ), .B(\U1/keyexpantion/SB0/n2372 ), .C(
        \U1/keyexpantion/SB0/n2371 ), .D(\U1/keyexpantion/SB0/n2370 ), .Y(
        \U1/keyexpantion/SB0/n2400 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U670  ( .A(\U1/keyexpantion/SB0/n2374 ), 
        .Y(\U1/keyexpantion/SB0/n2397 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U669  ( .A(\U1/keyexpantion/SB0/n2375 ), 
        .Y(\U1/keyexpantion/SB0/n2391 ) );
  OAI21B_X0P5M_A12TL \U1/keyexpantion/SB0/U668  ( .A0(
        \U1/keyexpantion/SB0/n2377 ), .A1(\U1/keyexpantion/SB0/n2514 ), .B0N(
        \U1/keyexpantion/SB0/n2376 ), .Y(\U1/keyexpantion/SB0/n2390 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U667  ( .A0(
        \U1/keyexpantion/SB0/n2521 ), .A1(\U1/keyexpantion/SB0/n2378 ), .B0(
        \U1/keyexpantion/SB0/n2428 ), .B1(\U1/keyexpantion/SB0/n2488 ), .C0(
        \U1/keyexpantion/SB0/n2502 ), .C1(\U1/keyexpantion/SB0/n2523 ), .Y(
        \U1/keyexpantion/SB0/n2389 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U666  ( .AN(
        \U1/keyexpantion/SB0/n2382 ), .B(\U1/keyexpantion/SB0/n2381 ), .C(
        \U1/keyexpantion/SB0/n2380 ), .D(\U1/keyexpantion/SB0/n2379 ), .Y(
        \U1/keyexpantion/SB0/n2388 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U665  ( .A(
        \U1/keyexpantion/SB0/n2386 ), .B(\U1/keyexpantion/SB0/n2385 ), .C(
        \U1/keyexpantion/SB0/n2384 ), .D(\U1/keyexpantion/SB0/n2383 ), .Y(
        \U1/keyexpantion/SB0/n2387 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U664  ( .A(\U1/keyexpantion/SB0/n2392 ), 
        .B(\U1/keyexpantion/SB0/n2391 ), .C(\U1/keyexpantion/SB0/n2390 ), .D(
        \U1/keyexpantion/SB0/n2389 ), .E(\U1/keyexpantion/SB0/n2388 ), .F(
        \U1/keyexpantion/SB0/n2387 ), .Y(\U1/keyexpantion/SB0/n2393 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U663  ( .A(\U1/keyexpantion/SB0/n2393 ), 
        .Y(\U1/keyexpantion/SB0/n2471 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U662  ( .A0(
        \U1/keyexpantion/SB0/n2461 ), .A1(\U1/keyexpantion/SB0/n2483 ), .B0(
        \U1/keyexpantion/SB0/n2523 ), .B1(\U1/keyexpantion/SB0/n2522 ), .Y(
        \U1/keyexpantion/SB0/n2394 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U661  ( .A0(
        \U1/keyexpantion/SB0/n2451 ), .A1(\U1/keyexpantion/SB0/n2395 ), .B0(
        \U1/keyexpantion/SB0/n2475 ), .B1(\U1/keyexpantion/SB0/n2497 ), .C0(
        \U1/keyexpantion/SB0/n2394 ), .Y(\U1/keyexpantion/SB0/n2396 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U660  ( .AN(
        \U1/keyexpantion/SB0/n2398 ), .B(\U1/keyexpantion/SB0/n2397 ), .C(
        \U1/keyexpantion/SB0/n2471 ), .D(\U1/keyexpantion/SB0/n2396 ), .Y(
        \U1/keyexpantion/SB0/n2399 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U659  ( .A(\U1/keyexpantion/SB0/n2404 ), 
        .B(\U1/keyexpantion/SB0/n2403 ), .C(\U1/keyexpantion/SB0/n2402 ), .D(
        \U1/keyexpantion/SB0/n2401 ), .E(\U1/keyexpantion/SB0/n2400 ), .F(
        \U1/keyexpantion/SB0/n2399 ), .Y(\U1/keyexpantion/SB0/n2469 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U658  ( .A(\U1/keyexpantion/SB0/n2405 ), 
        .Y(\U1/keyexpantion/SB0/n2409 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U657  ( .A0(
        \U1/keyexpantion/SB0/n2407 ), .A1(\U1/keyexpantion/SB0/n2406 ), .B0(
        \U1/keyexpantion/SB0/n2453 ), .B1(\U1/keyexpantion/SB0/n2412 ), .Y(
        \U1/keyexpantion/SB0/n2408 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U656  ( .A0(
        \U1/keyexpantion/SB0/n2502 ), .A1(\U1/keyexpantion/SB0/n2410 ), .B0(
        \U1/keyexpantion/SB0/n2409 ), .C0(\U1/keyexpantion/SB0/n2408 ), .Y(
        \U1/keyexpantion/SB0/n2424 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U655  ( .A0(
        \U1/keyexpantion/SB0/n2411 ), .A1(\U1/keyexpantion/SB0/n2474 ), .B0(
        \U1/keyexpantion/SB0/n2503 ), .Y(\U1/keyexpantion/SB0/n2416 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U654  ( .A0(
        \U1/keyexpantion/SB0/n2412 ), .A1(\U1/keyexpantion/SB0/n2477 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2415 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U653  ( .A(
        \U1/keyexpantion/SB0/n2416 ), .B(\U1/keyexpantion/SB0/n2415 ), .C(
        \U1/keyexpantion/SB0/n2414 ), .D(\U1/keyexpantion/SB0/n2413 ), .Y(
        \U1/keyexpantion/SB0/n2423 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U652  ( .A(\U1/keyexpantion/SB0/n2454 ), .B(\U1/keyexpantion/SB0/n2417 ), .Y(\U1/keyexpantion/SB0/n2421 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U651  ( .A(\U1/keyexpantion/SB0/n2418 ), .B(\U1/keyexpantion/SB0/n2459 ), .Y(\U1/keyexpantion/SB0/n2420 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U650  ( .A0(
        \U1/keyexpantion/SB0/n2421 ), .A1(\U1/keyexpantion/SB0/n2520 ), .B0(
        \U1/keyexpantion/SB0/n2420 ), .B1(\U1/keyexpantion/SB0/n2484 ), .C0(
        \U1/keyexpantion/SB0/n2419 ), .C1(\U1/keyexpantion/SB0/n2485 ), .Y(
        \U1/keyexpantion/SB0/n2422 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U649  ( .A(\U1/keyexpantion/SB0/n2493 ), 
        .B(\U1/keyexpantion/SB0/n2469 ), .C(\U1/keyexpantion/SB0/n2425 ), .D(
        \U1/keyexpantion/SB0/n2424 ), .E(\U1/keyexpantion/SB0/n2423 ), .F(
        \U1/keyexpantion/SB0/n2422 ), .Y(\U1/keyexpantion/ws [20]) );
  AOI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U648  ( .A1N(
        \U1/keyexpantion/SB0/n2427 ), .A0(\U1/keyexpantion/SB0/n2426 ), .B0(
        \U1/keyexpantion/SB0/n2483 ), .Y(\U1/keyexpantion/SB0/n2443 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U647  ( .A(\U1/keyexpantion/SB0/n2496 ), .B(\U1/keyexpantion/SB0/n2477 ), .Y(\U1/keyexpantion/SB0/n2430 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U646  ( .A0(
        \U1/keyexpantion/SB0/n2520 ), .A1(\U1/keyexpantion/SB0/n2431 ), .B0(
        \U1/keyexpantion/SB0/n2430 ), .B1(\U1/keyexpantion/SB0/n2523 ), .C0(
        \U1/keyexpantion/SB0/n2429 ), .C1(\U1/keyexpantion/SB0/n2428 ), .Y(
        \U1/keyexpantion/SB0/n2442 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U645  ( .A(\U1/keyexpantion/SB0/n2432 ), 
        .Y(\U1/keyexpantion/SB0/n2435 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U644  ( .AN(
        \U1/keyexpantion/SB0/n2436 ), .B(\U1/keyexpantion/SB0/n2435 ), .C(
        \U1/keyexpantion/SB0/n2434 ), .D(\U1/keyexpantion/SB0/n2433 ), .Y(
        \U1/keyexpantion/SB0/n2441 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U643  ( .A(
        \U1/keyexpantion/SB0/n2439 ), .B(\U1/keyexpantion/SB0/n2438 ), .C(
        \U1/keyexpantion/SB0/n2437 ), .Y(\U1/keyexpantion/SB0/n2440 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U642  ( .A(\U1/keyexpantion/SB0/n2445 ), 
        .B(\U1/keyexpantion/SB0/n2444 ), .C(\U1/keyexpantion/SB0/n2443 ), .D(
        \U1/keyexpantion/SB0/n2442 ), .E(\U1/keyexpantion/SB0/n2441 ), .F(
        \U1/keyexpantion/SB0/n2440 ), .Y(\U1/keyexpantion/SB0/n2494 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U641  ( .A(\U1/keyexpantion/SB0/n2446 ), 
        .Y(\U1/keyexpantion/SB0/n2448 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U640  ( .A0(
        \U1/keyexpantion/SB0/n2507 ), .A1(\U1/keyexpantion/SB0/n2504 ), .B0(
        \U1/keyexpantion/SB0/n2508 ), .B1(\U1/keyexpantion/SB0/n2506 ), .Y(
        \U1/keyexpantion/SB0/n2447 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U639  ( .A0(
        \U1/keyexpantion/SB0/n2483 ), .A1(\U1/keyexpantion/SB0/n2449 ), .B0(
        \U1/keyexpantion/SB0/n2448 ), .C0(\U1/keyexpantion/SB0/n2447 ), .Y(
        \U1/keyexpantion/SB0/n2468 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U638  ( .A0(
        \U1/keyexpantion/SB0/n2451 ), .A1(\U1/keyexpantion/SB0/n2507 ), .B0(
        \U1/keyexpantion/SB0/n2450 ), .Y(\U1/keyexpantion/SB0/n2457 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U637  ( .A0(
        \U1/keyexpantion/SB0/n2454 ), .A1(\U1/keyexpantion/SB0/n2453 ), .B0(
        \U1/keyexpantion/SB0/n2452 ), .Y(\U1/keyexpantion/SB0/n2456 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U636  ( .AN(
        \U1/keyexpantion/SB0/n2458 ), .B(\U1/keyexpantion/SB0/n2457 ), .C(
        \U1/keyexpantion/SB0/n2456 ), .D(\U1/keyexpantion/SB0/n2455 ), .Y(
        \U1/keyexpantion/SB0/n2467 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U635  ( .A0(
        \U1/keyexpantion/SB0/n2503 ), .A1(\U1/keyexpantion/SB0/n2460 ), .B0(
        \U1/keyexpantion/SB0/n2459 ), .Y(\U1/keyexpantion/SB0/n2464 ) );
  OA22_X0P5M_A12TL \U1/keyexpantion/SB0/U634  ( .A0(
        \U1/keyexpantion/SB0/n2485 ), .A1(\U1/keyexpantion/SB0/n2462 ), .B0(
        \U1/keyexpantion/SB0/n2522 ), .B1(\U1/keyexpantion/SB0/n2461 ), .Y(
        \U1/keyexpantion/SB0/n2463 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U633  ( .A0(
        \U1/keyexpantion/SB0/n2465 ), .A1(\U1/keyexpantion/SB0/n2484 ), .B0(
        \U1/keyexpantion/SB0/n2464 ), .C0(\U1/keyexpantion/SB0/n2463 ), .Y(
        \U1/keyexpantion/SB0/n2466 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U632  ( .A(\U1/keyexpantion/SB0/n2494 ), 
        .B(\U1/keyexpantion/SB0/n2470 ), .C(\U1/keyexpantion/SB0/n2469 ), .D(
        \U1/keyexpantion/SB0/n2468 ), .E(\U1/keyexpantion/SB0/n2467 ), .F(
        \U1/keyexpantion/SB0/n2466 ), .Y(\U1/keyexpantion/ws [21]) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U631  ( .A0(
        \U1/keyexpantion/SB0/n2473 ), .A1(\U1/keyexpantion/SB0/n2513 ), .B0(
        \U1/keyexpantion/SB0/n2472 ), .B1(\U1/keyexpantion/SB0/n2520 ), .C0(
        \U1/keyexpantion/SB0/n2471 ), .Y(\U1/keyexpantion/SB0/n2491 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U630  ( .A0(
        \U1/keyexpantion/SB0/n2474 ), .A1(\U1/keyexpantion/SB0/n2518 ), .B0(
        \U1/keyexpantion/SB0/n2507 ), .Y(\U1/keyexpantion/SB0/n2482 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U629  ( .A0(
        \U1/keyexpantion/SB0/n2498 ), .A1(\U1/keyexpantion/SB0/n2475 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2481 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U628  ( .A0(
        \U1/keyexpantion/SB0/n2478 ), .A1(\U1/keyexpantion/SB0/n2477 ), .B0(
        \U1/keyexpantion/SB0/n2476 ), .Y(\U1/keyexpantion/SB0/n2480 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U627  ( .A(
        \U1/keyexpantion/SB0/n2482 ), .B(\U1/keyexpantion/SB0/n2481 ), .C(
        \U1/keyexpantion/SB0/n2480 ), .D(\U1/keyexpantion/SB0/n2479 ), .Y(
        \U1/keyexpantion/SB0/n2490 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U626  ( .A(
        \U1/keyexpantion/SB0/n2513 ), .B(\U1/keyexpantion/SB0/n2483 ), .Y(
        \U1/keyexpantion/SB0/n2515 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U625  ( .A(\U1/keyexpantion/SB0/n2503 ), .B(\U1/keyexpantion/SB0/n2515 ), .Y(\U1/keyexpantion/SB0/n2487 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U624  ( .A0(
        \U1/keyexpantion/SB0/n2501 ), .A1(\U1/keyexpantion/SB0/n2488 ), .B0(
        \U1/keyexpantion/SB0/n2487 ), .B1(\U1/keyexpantion/SB0/n2486 ), .C0(
        \U1/keyexpantion/SB0/n2485 ), .C1(\U1/keyexpantion/SB0/n2484 ), .Y(
        \U1/keyexpantion/SB0/n2489 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U623  ( .A(\U1/keyexpantion/SB0/n2494 ), 
        .B(\U1/keyexpantion/SB0/n2493 ), .C(\U1/keyexpantion/SB0/n2492 ), .D(
        \U1/keyexpantion/SB0/n2491 ), .E(\U1/keyexpantion/SB0/n2490 ), .F(
        \U1/keyexpantion/SB0/n2489 ), .Y(\U1/keyexpantion/ws [22]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U622  ( .A0(
        \U1/keyexpantion/SB0/n2498 ), .A1(\U1/keyexpantion/SB0/n2497 ), .B0(
        \U1/keyexpantion/SB0/n2496 ), .B1(\U1/keyexpantion/SB0/n2495 ), .Y(
        \U1/keyexpantion/SB0/n2499 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U621  ( .A0(
        \U1/keyexpantion/SB0/n2502 ), .A1(\U1/keyexpantion/SB0/n2501 ), .B0(
        \U1/keyexpantion/SB0/n2500 ), .C0(\U1/keyexpantion/SB0/n2499 ), .Y(
        \U1/keyexpantion/SB0/n2526 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U620  ( .A1N(
        \U1/keyexpantion/SB0/n2505 ), .A0(\U1/keyexpantion/SB0/n2504 ), .B0(
        \U1/keyexpantion/SB0/n2503 ), .Y(\U1/keyexpantion/SB0/n2512 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U619  ( .A0(
        \U1/keyexpantion/SB0/n2508 ), .A1(\U1/keyexpantion/SB0/n2507 ), .B0(
        \U1/keyexpantion/SB0/n2506 ), .Y(\U1/keyexpantion/SB0/n2511 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U618  ( .A(
        \U1/keyexpantion/SB0/n2512 ), .B(\U1/keyexpantion/SB0/n2511 ), .C(
        \U1/keyexpantion/SB0/n2510 ), .D(\U1/keyexpantion/SB0/n2509 ), .Y(
        \U1/keyexpantion/SB0/n2525 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U617  ( .A(
        \U1/keyexpantion/SB0/n2514 ), .B(\U1/keyexpantion/SB0/n2513 ), .Y(
        \U1/keyexpantion/SB0/n2517 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U616  ( .A0(
        \U1/keyexpantion/SB0/n2518 ), .A1(\U1/keyexpantion/SB0/n2517 ), .B0(
        \U1/keyexpantion/SB0/n2516 ), .B1(\U1/keyexpantion/SB0/n2515 ), .Y(
        \U1/keyexpantion/SB0/n2519 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U615  ( .A0(
        \U1/keyexpantion/SB0/n2523 ), .A1(\U1/keyexpantion/SB0/n2522 ), .B0(
        \U1/keyexpantion/SB0/n2521 ), .B1(\U1/keyexpantion/SB0/n2520 ), .C0(
        \U1/keyexpantion/SB0/n2519 ), .Y(\U1/keyexpantion/SB0/n2524 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U614  ( .A(\U1/keyexpantion/SB0/n2529 ), 
        .B(\U1/keyexpantion/SB0/n2528 ), .C(\U1/keyexpantion/SB0/n2527 ), .D(
        \U1/keyexpantion/SB0/n2526 ), .E(\U1/keyexpantion/SB0/n2525 ), .F(
        \U1/keyexpantion/SB0/n2524 ), .Y(\U1/keyexpantion/ws [23]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U613  ( .A(\U1/rkey [23]), .B(
        \U1/rkey [22]), .Y(\U1/keyexpantion/SB0/n2548 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U612  ( .A(\U1/rkey [21]), .B(
        \U1/rkey [20]), .Y(\U1/keyexpantion/SB0/n2539 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U611  ( .A(
        \U1/keyexpantion/SB0/n2548 ), .B(\U1/keyexpantion/SB0/n2539 ), .Y(
        \U1/keyexpantion/SB0/n2613 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U610  ( .A(\U1/rkey [17]), .Y(
        \U1/keyexpantion/SB0/n2533 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U609  ( .A(\U1/rkey [16]), .Y(
        \U1/keyexpantion/SB0/n2530 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U608  ( .A(\U1/keyexpantion/SB0/n2533 ), .B(\U1/keyexpantion/SB0/n2530 ), .Y(\U1/keyexpantion/SB0/n2540 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U607  ( .A(\U1/rkey [19]), .B(
        \U1/rkey [18]), .Y(\U1/keyexpantion/SB0/n2560 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U606  ( .A(
        \U1/keyexpantion/SB0/n2540 ), .B(\U1/keyexpantion/SB0/n2560 ), .Y(
        \U1/keyexpantion/SB0/n2916 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U605  ( .A(\U1/keyexpantion/SB0/n2613 ), .B(\U1/keyexpantion/SB0/n2916 ), .Y(\U1/keyexpantion/SB0/n2702 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U604  ( .A(\U1/rkey [18]), .B(
        \U1/rkey [19]), .Y(\U1/keyexpantion/SB0/n2543 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U603  ( .A(
        \U1/keyexpantion/SB0/n2543 ), .B(\U1/keyexpantion/SB0/n2540 ), .Y(
        \U1/keyexpantion/SB0/n2833 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U602  ( .A(\U1/rkey [23]), .Y(
        \U1/keyexpantion/SB0/n2536 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U601  ( .A(\U1/keyexpantion/SB0/n2536 ), .B(\U1/rkey [22]), .Y(\U1/keyexpantion/SB0/n2566 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U600  ( .A(
        \U1/keyexpantion/SB0/n2566 ), .B(\U1/keyexpantion/SB0/n2539 ), .Y(
        \U1/keyexpantion/SB0/n2612 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U599  ( .A(\U1/keyexpantion/SB0/n2833 ), .B(\U1/keyexpantion/SB0/n2612 ), .Y(\U1/keyexpantion/SB0/n2799 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U598  ( .A(\U1/rkey [19]), .Y(
        \U1/keyexpantion/SB0/n2531 ) );
  AND2_X0P5M_A12TL \U1/keyexpantion/SB0/U597  ( .A(\U1/rkey [18]), .B(
        \U1/keyexpantion/SB0/n2531 ), .Y(\U1/keyexpantion/SB0/n2541 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U596  ( .A(
        \U1/keyexpantion/SB0/n2540 ), .B(\U1/keyexpantion/SB0/n2541 ), .Y(
        \U1/keyexpantion/SB0/n2764 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U595  ( .A(\U1/keyexpantion/SB0/n2764 ), 
        .Y(\U1/keyexpantion/SB0/n2950 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U594  ( .A(\U1/rkey [20]), .Y(
        \U1/keyexpantion/SB0/n2532 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U593  ( .A(\U1/keyexpantion/SB0/n2532 ), .B(\U1/rkey [21]), .Y(\U1/keyexpantion/SB0/n2547 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U592  ( .A(\U1/rkey [22]), .Y(
        \U1/keyexpantion/SB0/n2535 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U591  ( .A(\U1/keyexpantion/SB0/n2535 ), .B(\U1/rkey [23]), .Y(\U1/keyexpantion/SB0/n2557 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U590  ( .A(
        \U1/keyexpantion/SB0/n2547 ), .B(\U1/keyexpantion/SB0/n2557 ), .Y(
        \U1/keyexpantion/SB0/n2785 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U589  ( .A(\U1/keyexpantion/SB0/n2785 ), 
        .Y(\U1/keyexpantion/SB0/n2883 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U588  ( .A(
        \U1/keyexpantion/SB0/n2950 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2742 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U587  ( .A(\U1/keyexpantion/SB0/n2613 ), 
        .Y(\U1/keyexpantion/SB0/n2919 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U586  ( .A(\U1/rkey [17]), .B(
        \U1/rkey [16]), .Y(\U1/keyexpantion/SB0/n2544 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U585  ( .A(
        \U1/keyexpantion/SB0/n2544 ), .B(\U1/keyexpantion/SB0/n2560 ), .Y(
        \U1/keyexpantion/SB0/n2851 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U584  ( .A(\U1/keyexpantion/SB0/n2851 ), 
        .Y(\U1/keyexpantion/SB0/n2960 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U583  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2960 ), .Y(
        \U1/keyexpantion/SB0/n2856 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U582  ( .A(\U1/keyexpantion/SB0/n2530 ), .B(\U1/rkey [17]), .Y(\U1/keyexpantion/SB0/n2559 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U581  ( .A(
        \U1/keyexpantion/SB0/n2541 ), .B(\U1/keyexpantion/SB0/n2559 ), .Y(
        \U1/keyexpantion/SB0/n2751 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U580  ( .A(\U1/keyexpantion/SB0/n2751 ), 
        .Y(\U1/keyexpantion/SB0/n2840 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U579  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2720 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U578  ( .A(
        \U1/keyexpantion/SB0/n2742 ), .B(\U1/keyexpantion/SB0/n2856 ), .C(
        \U1/keyexpantion/SB0/n2720 ), .Y(\U1/keyexpantion/SB0/n2579 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U577  ( .A(
        \U1/keyexpantion/SB0/n2539 ), .B(\U1/keyexpantion/SB0/n2557 ), .Y(
        \U1/keyexpantion/SB0/n2784 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U576  ( .A(\U1/keyexpantion/SB0/n2531 ), .B(\U1/rkey [18]), .Y(\U1/keyexpantion/SB0/n2550 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U575  ( .A(
        \U1/keyexpantion/SB0/n2550 ), .B(\U1/keyexpantion/SB0/n2559 ), .Y(
        \U1/keyexpantion/SB0/n2782 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U574  ( .A(\U1/keyexpantion/SB0/n2784 ), .B(\U1/keyexpantion/SB0/n2782 ), .Y(\U1/keyexpantion/SB0/n2697 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U573  ( .A(\U1/keyexpantion/SB0/n2612 ), 
        .Y(\U1/keyexpantion/SB0/n2921 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U572  ( .A(\U1/rkey [21]), .Y(
        \U1/keyexpantion/SB0/n2534 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U571  ( .A(\U1/keyexpantion/SB0/n2532 ), .B(\U1/keyexpantion/SB0/n2534 ), .Y(\U1/keyexpantion/SB0/n2558 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U570  ( .A(
        \U1/keyexpantion/SB0/n2548 ), .B(\U1/keyexpantion/SB0/n2558 ), .Y(
        \U1/keyexpantion/SB0/n2964 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U569  ( .A(\U1/keyexpantion/SB0/n2964 ), 
        .Y(\U1/keyexpantion/SB0/n2874 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U568  ( .A(\U1/keyexpantion/SB0/n2533 ), .B(\U1/rkey [16]), .Y(\U1/keyexpantion/SB0/n2549 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U567  ( .A(
        \U1/keyexpantion/SB0/n2549 ), .B(\U1/keyexpantion/SB0/n2560 ), .Y(
        \U1/keyexpantion/SB0/n2929 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U566  ( .A(\U1/keyexpantion/SB0/n2929 ), 
        .Y(\U1/keyexpantion/SB0/n2756 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U565  ( .A0(
        \U1/keyexpantion/SB0/n2921 ), .A1(\U1/keyexpantion/SB0/n2874 ), .B0(
        \U1/keyexpantion/SB0/n2756 ), .Y(\U1/keyexpantion/SB0/n2538 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U564  ( .A(
        \U1/keyexpantion/SB0/n2544 ), .B(\U1/keyexpantion/SB0/n2541 ), .Y(
        \U1/keyexpantion/SB0/n2917 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U563  ( .A(\U1/keyexpantion/SB0/n2917 ), 
        .Y(\U1/keyexpantion/SB0/n2882 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U562  ( .A(\U1/keyexpantion/SB0/n2534 ), .B(\U1/rkey [20]), .Y(\U1/keyexpantion/SB0/n2565 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U561  ( .A(
        \U1/keyexpantion/SB0/n2557 ), .B(\U1/keyexpantion/SB0/n2565 ), .Y(
        \U1/keyexpantion/SB0/n2957 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U560  ( .A(
        \U1/keyexpantion/SB0/n2784 ), .B(\U1/keyexpantion/SB0/n2957 ), .Y(
        \U1/keyexpantion/SB0/n2675 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U559  ( .A(\U1/keyexpantion/SB0/n2536 ), .B(\U1/keyexpantion/SB0/n2535 ), .Y(\U1/keyexpantion/SB0/n2556 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U558  ( .A(
        \U1/keyexpantion/SB0/n2547 ), .B(\U1/keyexpantion/SB0/n2556 ), .Y(
        \U1/keyexpantion/SB0/n2932 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U557  ( .A(\U1/keyexpantion/SB0/n2932 ), 
        .Y(\U1/keyexpantion/SB0/n2656 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U556  ( .A0(
        \U1/keyexpantion/SB0/n2882 ), .A1(\U1/keyexpantion/SB0/n2675 ), .B0(
        \U1/keyexpantion/SB0/n2656 ), .B1(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2537 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U555  ( .AN(
        \U1/keyexpantion/SB0/n2697 ), .B(\U1/keyexpantion/SB0/n2538 ), .C(
        \U1/keyexpantion/SB0/n2537 ), .Y(\U1/keyexpantion/SB0/n2578 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U554  ( .A(
        \U1/keyexpantion/SB0/n2539 ), .B(\U1/keyexpantion/SB0/n2556 ), .Y(
        \U1/keyexpantion/SB0/n2801 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U553  ( .A(
        \U1/keyexpantion/SB0/n2543 ), .B(\U1/keyexpantion/SB0/n2544 ), .Y(
        \U1/keyexpantion/SB0/n2967 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U552  ( .A(
        \U1/keyexpantion/SB0/n2566 ), .B(\U1/keyexpantion/SB0/n2547 ), .Y(
        \U1/keyexpantion/SB0/n2852 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U551  ( .A(
        \U1/keyexpantion/SB0/n2543 ), .B(\U1/keyexpantion/SB0/n2549 ), .Y(
        \U1/keyexpantion/SB0/n2849 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U550  ( .A(
        \U1/keyexpantion/SB0/n2540 ), .B(\U1/keyexpantion/SB0/n2550 ), .Y(
        \U1/keyexpantion/SB0/n2854 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U549  ( .A(\U1/keyexpantion/SB0/n2854 ), 
        .Y(\U1/keyexpantion/SB0/n2834 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U548  ( .A(\U1/keyexpantion/SB0/n2957 ), 
        .Y(\U1/keyexpantion/SB0/n2670 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U547  ( .A(
        \U1/keyexpantion/SB0/n2541 ), .B(\U1/keyexpantion/SB0/n2549 ), .Y(
        \U1/keyexpantion/SB0/n2872 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U546  ( .A(\U1/keyexpantion/SB0/n2872 ), 
        .Y(\U1/keyexpantion/SB0/n2918 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U545  ( .A0(
        \U1/keyexpantion/SB0/n2834 ), .A1(\U1/keyexpantion/SB0/n2919 ), .B0(
        \U1/keyexpantion/SB0/n2670 ), .B1(\U1/keyexpantion/SB0/n2918 ), .Y(
        \U1/keyexpantion/SB0/n2542 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U544  ( .A0(
        \U1/keyexpantion/SB0/n2801 ), .A1(\U1/keyexpantion/SB0/n2967 ), .B0(
        \U1/keyexpantion/SB0/n2852 ), .B1(\U1/keyexpantion/SB0/n2849 ), .C0(
        \U1/keyexpantion/SB0/n2542 ), .Y(\U1/keyexpantion/SB0/n2577 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U543  ( .A(\U1/keyexpantion/SB0/n2854 ), .B(\U1/keyexpantion/SB0/n2801 ), .Y(\U1/keyexpantion/SB0/n2663 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U542  ( .A(\U1/keyexpantion/SB0/n2849 ), .B(\U1/keyexpantion/SB0/n2784 ), .Y(\U1/keyexpantion/SB0/n2673 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U541  ( .A(\U1/keyexpantion/SB0/n2673 ), 
        .Y(\U1/keyexpantion/SB0/n2546 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U540  ( .A(
        \U1/keyexpantion/SB0/n2543 ), .B(\U1/keyexpantion/SB0/n2559 ), .Y(
        \U1/keyexpantion/SB0/n2945 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U539  ( .A(\U1/keyexpantion/SB0/n2945 ), 
        .Y(\U1/keyexpantion/SB0/n2873 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U538  ( .A(
        \U1/keyexpantion/SB0/n2544 ), .B(\U1/keyexpantion/SB0/n2550 ), .Y(
        \U1/keyexpantion/SB0/n2930 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U537  ( .A(\U1/keyexpantion/SB0/n2930 ), 
        .Y(\U1/keyexpantion/SB0/n2941 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U536  ( .A0(
        \U1/keyexpantion/SB0/n2873 ), .A1(\U1/keyexpantion/SB0/n2941 ), .B0(
        \U1/keyexpantion/SB0/n2874 ), .Y(\U1/keyexpantion/SB0/n2545 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U535  ( .A(
        \U1/keyexpantion/SB0/n2548 ), .B(\U1/keyexpantion/SB0/n2565 ), .Y(
        \U1/keyexpantion/SB0/n2946 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U534  ( .A(\U1/keyexpantion/SB0/n2946 ), 
        .Y(\U1/keyexpantion/SB0/n2875 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U533  ( .A(
        \U1/keyexpantion/SB0/n2875 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2690 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U532  ( .AN(
        \U1/keyexpantion/SB0/n2663 ), .B(\U1/keyexpantion/SB0/n2546 ), .C(
        \U1/keyexpantion/SB0/n2545 ), .D(\U1/keyexpantion/SB0/n2690 ), .Y(
        \U1/keyexpantion/SB0/n2555 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U531  ( .A(
        \U1/keyexpantion/SB0/n2558 ), .B(\U1/keyexpantion/SB0/n2556 ), .Y(
        \U1/keyexpantion/SB0/n2966 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U530  ( .A(
        \U1/keyexpantion/SB0/n2548 ), .B(\U1/keyexpantion/SB0/n2547 ), .Y(
        \U1/keyexpantion/SB0/n2958 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U529  ( .A0(
        \U1/keyexpantion/SB0/n2612 ), .A1(\U1/keyexpantion/SB0/n2764 ), .B0(
        \U1/keyexpantion/SB0/n2966 ), .B1(\U1/keyexpantion/SB0/n2854 ), .C0(
        \U1/keyexpantion/SB0/n2958 ), .C1(\U1/keyexpantion/SB0/n2872 ), .Y(
        \U1/keyexpantion/SB0/n2554 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U528  ( .A(\U1/keyexpantion/SB0/n2917 ), .B(\U1/keyexpantion/SB0/n2612 ), .Y(\U1/keyexpantion/SB0/n2748 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U527  ( .A(
        \U1/keyexpantion/SB0/n2670 ), .B(\U1/keyexpantion/SB0/n2834 ), .Y(
        \U1/keyexpantion/SB0/n2701 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U526  ( .A(
        \U1/keyexpantion/SB0/n2918 ), .B(\U1/keyexpantion/SB0/n2919 ), .Y(
        \U1/keyexpantion/SB0/n2721 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U525  ( .A(\U1/keyexpantion/SB0/n2852 ), 
        .Y(\U1/keyexpantion/SB0/n2947 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U524  ( .A(
        \U1/keyexpantion/SB0/n2947 ), .B(\U1/keyexpantion/SB0/n2756 ), .Y(
        \U1/keyexpantion/SB0/n2759 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U523  ( .AN(
        \U1/keyexpantion/SB0/n2748 ), .B(\U1/keyexpantion/SB0/n2701 ), .C(
        \U1/keyexpantion/SB0/n2721 ), .D(\U1/keyexpantion/SB0/n2759 ), .Y(
        \U1/keyexpantion/SB0/n2553 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U522  ( .A(
        \U1/keyexpantion/SB0/n2566 ), .B(\U1/keyexpantion/SB0/n2558 ), .Y(
        \U1/keyexpantion/SB0/n2671 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U521  ( .A(\U1/keyexpantion/SB0/n2671 ), .B(\U1/keyexpantion/SB0/n2929 ), .Y(\U1/keyexpantion/SB0/n2825 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U520  ( .A(
        \U1/keyexpantion/SB0/n2550 ), .B(\U1/keyexpantion/SB0/n2549 ), .Y(
        \U1/keyexpantion/SB0/n2965 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U519  ( .A(\U1/keyexpantion/SB0/n2932 ), .B(\U1/keyexpantion/SB0/n2965 ), .Y(\U1/keyexpantion/SB0/n2790 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U518  ( .A(\U1/keyexpantion/SB0/n2790 ), 
        .Y(\U1/keyexpantion/SB0/n2551 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U517  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2756 ), .Y(
        \U1/keyexpantion/SB0/n2809 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U516  ( .A(\U1/keyexpantion/SB0/n2965 ), 
        .Y(\U1/keyexpantion/SB0/n2948 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U515  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2948 ), .Y(
        \U1/keyexpantion/SB0/n2860 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U514  ( .AN(
        \U1/keyexpantion/SB0/n2825 ), .B(\U1/keyexpantion/SB0/n2551 ), .C(
        \U1/keyexpantion/SB0/n2809 ), .D(\U1/keyexpantion/SB0/n2860 ), .Y(
        \U1/keyexpantion/SB0/n2552 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U513  ( .A(\U1/keyexpantion/SB0/n2555 ), 
        .B(\U1/keyexpantion/SB0/n2554 ), .C(\U1/keyexpantion/SB0/n2553 ), .D(
        \U1/keyexpantion/SB0/n2552 ), .Y(\U1/keyexpantion/SB0/n2652 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U512  ( .A(\U1/keyexpantion/SB0/n2851 ), .B(\U1/keyexpantion/SB0/n2671 ), .Y(\U1/keyexpantion/SB0/n2859 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U511  ( .A(
        \U1/keyexpantion/SB0/n2565 ), .B(\U1/keyexpantion/SB0/n2556 ), .Y(
        \U1/keyexpantion/SB0/n2767 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U510  ( .A(\U1/keyexpantion/SB0/n2833 ), .B(\U1/keyexpantion/SB0/n2767 ), .Y(\U1/keyexpantion/SB0/n2738 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U509  ( .A(\U1/keyexpantion/SB0/n2966 ), 
        .Y(\U1/keyexpantion/SB0/n2922 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U508  ( .A(
        \U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2882 ), .Y(
        \U1/keyexpantion/SB0/n2687 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U507  ( .A0(
        \U1/keyexpantion/SB0/n2767 ), .A1(\U1/keyexpantion/SB0/n2965 ), .B0(
        \U1/keyexpantion/SB0/n2687 ), .Y(\U1/keyexpantion/SB0/n2564 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U506  ( .A(\U1/keyexpantion/SB0/n2782 ), 
        .Y(\U1/keyexpantion/SB0/n2877 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U505  ( .A(
        \U1/keyexpantion/SB0/n2877 ), .B(\U1/keyexpantion/SB0/n2921 ), .Y(
        \U1/keyexpantion/SB0/n2878 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U504  ( .A(
        \U1/keyexpantion/SB0/n2921 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2837 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U503  ( .A(
        \U1/keyexpantion/SB0/n2558 ), .B(\U1/keyexpantion/SB0/n2557 ), .Y(
        \U1/keyexpantion/SB0/n2928 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U502  ( .A(\U1/keyexpantion/SB0/n2928 ), 
        .Y(\U1/keyexpantion/SB0/n2682 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U501  ( .A(
        \U1/keyexpantion/SB0/n2873 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2706 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U500  ( .A(\U1/keyexpantion/SB0/n2916 ), 
        .Y(\U1/keyexpantion/SB0/n2876 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U499  ( .A(
        \U1/keyexpantion/SB0/n2876 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2770 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U498  ( .A(
        \U1/keyexpantion/SB0/n2878 ), .B(\U1/keyexpantion/SB0/n2837 ), .C(
        \U1/keyexpantion/SB0/n2706 ), .D(\U1/keyexpantion/SB0/n2770 ), .Y(
        \U1/keyexpantion/SB0/n2563 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U497  ( .A(
        \U1/keyexpantion/SB0/n2918 ), .B(\U1/keyexpantion/SB0/n2875 ), .Y(
        \U1/keyexpantion/SB0/n2804 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U496  ( .A(
        \U1/keyexpantion/SB0/n2960 ), .B(\U1/keyexpantion/SB0/n2875 ), .Y(
        \U1/keyexpantion/SB0/n2795 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U495  ( .A(\U1/keyexpantion/SB0/n2958 ), 
        .Y(\U1/keyexpantion/SB0/n2951 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U494  ( .A(
        \U1/keyexpantion/SB0/n2834 ), .B(\U1/keyexpantion/SB0/n2951 ), .Y(
        \U1/keyexpantion/SB0/n2667 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U493  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2873 ), .Y(
        \U1/keyexpantion/SB0/n2778 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U492  ( .A(
        \U1/keyexpantion/SB0/n2804 ), .B(\U1/keyexpantion/SB0/n2795 ), .C(
        \U1/keyexpantion/SB0/n2667 ), .D(\U1/keyexpantion/SB0/n2778 ), .Y(
        \U1/keyexpantion/SB0/n2562 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U491  ( .A(\U1/keyexpantion/SB0/n2849 ), 
        .Y(\U1/keyexpantion/SB0/n2818 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U490  ( .A(
        \U1/keyexpantion/SB0/n2670 ), .B(\U1/keyexpantion/SB0/n2818 ), .Y(
        \U1/keyexpantion/SB0/n2654 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U489  ( .A(
        \U1/keyexpantion/SB0/n2560 ), .B(\U1/keyexpantion/SB0/n2559 ), .Y(
        \U1/keyexpantion/SB0/n2884 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U488  ( .A(\U1/keyexpantion/SB0/n2884 ), 
        .Y(\U1/keyexpantion/SB0/n2939 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U487  ( .A(
        \U1/keyexpantion/SB0/n2670 ), .B(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2718 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U486  ( .A(\U1/keyexpantion/SB0/n2833 ), 
        .Y(\U1/keyexpantion/SB0/n2962 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U485  ( .A(
        \U1/keyexpantion/SB0/n2962 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2753 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U484  ( .A(
        \U1/keyexpantion/SB0/n2874 ), .B(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2923 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U483  ( .A(
        \U1/keyexpantion/SB0/n2654 ), .B(\U1/keyexpantion/SB0/n2718 ), .C(
        \U1/keyexpantion/SB0/n2753 ), .D(\U1/keyexpantion/SB0/n2923 ), .Y(
        \U1/keyexpantion/SB0/n2561 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U482  ( .A(\U1/keyexpantion/SB0/n2859 ), 
        .B(\U1/keyexpantion/SB0/n2738 ), .C(\U1/keyexpantion/SB0/n2564 ), .D(
        \U1/keyexpantion/SB0/n2563 ), .E(\U1/keyexpantion/SB0/n2562 ), .F(
        \U1/keyexpantion/SB0/n2561 ), .Y(\U1/keyexpantion/SB0/n2641 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U481  ( .A(\U1/keyexpantion/SB0/n2641 ), 
        .Y(\U1/keyexpantion/SB0/n2575 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U480  ( .A(\U1/keyexpantion/SB0/n2930 ), .B(\U1/keyexpantion/SB0/n2767 ), .Y(\U1/keyexpantion/SB0/n2664 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U479  ( .A(
        \U1/keyexpantion/SB0/n2566 ), .B(\U1/keyexpantion/SB0/n2565 ), .Y(
        \U1/keyexpantion/SB0/n2927 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U478  ( .A(\U1/keyexpantion/SB0/n2927 ), .B(\U1/keyexpantion/SB0/n2782 ), .Y(\U1/keyexpantion/SB0/n2791 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U477  ( .A(\U1/keyexpantion/SB0/n2791 ), 
        .Y(\U1/keyexpantion/SB0/n2568 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U476  ( .A(\U1/keyexpantion/SB0/n2784 ), 
        .Y(\U1/keyexpantion/SB0/n2952 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U475  ( .A0(
        \U1/keyexpantion/SB0/n2682 ), .A1(\U1/keyexpantion/SB0/n2952 ), .B0(
        \U1/keyexpantion/SB0/n2939 ), .Y(\U1/keyexpantion/SB0/n2567 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U474  ( .A(
        \U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2818 ), .Y(
        \U1/keyexpantion/SB0/n2689 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U473  ( .AN(
        \U1/keyexpantion/SB0/n2664 ), .B(\U1/keyexpantion/SB0/n2568 ), .C(
        \U1/keyexpantion/SB0/n2567 ), .D(\U1/keyexpantion/SB0/n2689 ), .Y(
        \U1/keyexpantion/SB0/n2572 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U472  ( .A0(
        \U1/keyexpantion/SB0/n2916 ), .A1(\U1/keyexpantion/SB0/n2964 ), .B0(
        \U1/keyexpantion/SB0/n2801 ), .B1(\U1/keyexpantion/SB0/n2849 ), .C0(
        \U1/keyexpantion/SB0/n2929 ), .C1(\U1/keyexpantion/SB0/n2946 ), .Y(
        \U1/keyexpantion/SB0/n2571 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U471  ( .A(\U1/keyexpantion/SB0/n2964 ), .B(\U1/keyexpantion/SB0/n2967 ), .Y(\U1/keyexpantion/SB0/n2729 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U470  ( .A(
        \U1/keyexpantion/SB0/n2952 ), .B(\U1/keyexpantion/SB0/n2873 ), .Y(
        \U1/keyexpantion/SB0/n2862 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U469  ( .A(
        \U1/keyexpantion/SB0/n2834 ), .B(\U1/keyexpantion/SB0/n2952 ), .Y(
        \U1/keyexpantion/SB0/n2796 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U468  ( .A(
        \U1/keyexpantion/SB0/n2818 ), .B(\U1/keyexpantion/SB0/n2919 ), .Y(
        \U1/keyexpantion/SB0/n2668 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U467  ( .AN(
        \U1/keyexpantion/SB0/n2729 ), .B(\U1/keyexpantion/SB0/n2862 ), .C(
        \U1/keyexpantion/SB0/n2796 ), .D(\U1/keyexpantion/SB0/n2668 ), .Y(
        \U1/keyexpantion/SB0/n2570 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U466  ( .A(
        \U1/keyexpantion/SB0/n2962 ), .B(\U1/keyexpantion/SB0/n2947 ), .Y(
        \U1/keyexpantion/SB0/n2741 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U465  ( .A(
        \U1/keyexpantion/SB0/n2818 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2808 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U464  ( .A(
        \U1/keyexpantion/SB0/n2670 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2709 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U463  ( .A(
        \U1/keyexpantion/SB0/n2877 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2754 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U462  ( .A(
        \U1/keyexpantion/SB0/n2741 ), .B(\U1/keyexpantion/SB0/n2808 ), .C(
        \U1/keyexpantion/SB0/n2709 ), .D(\U1/keyexpantion/SB0/n2754 ), .Y(
        \U1/keyexpantion/SB0/n2569 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U461  ( .A(\U1/keyexpantion/SB0/n2572 ), 
        .B(\U1/keyexpantion/SB0/n2571 ), .C(\U1/keyexpantion/SB0/n2570 ), .D(
        \U1/keyexpantion/SB0/n2569 ), .Y(\U1/keyexpantion/SB0/n2573 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U460  ( .A(\U1/keyexpantion/SB0/n2573 ), 
        .Y(\U1/keyexpantion/SB0/n2944 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U459  ( .A(
        \U1/keyexpantion/SB0/n2960 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2574 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U458  ( .AN(
        \U1/keyexpantion/SB0/n2652 ), .B(\U1/keyexpantion/SB0/n2575 ), .C(
        \U1/keyexpantion/SB0/n2944 ), .D(\U1/keyexpantion/SB0/n2574 ), .Y(
        \U1/keyexpantion/SB0/n2576 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U457  ( .A(\U1/keyexpantion/SB0/n2702 ), 
        .B(\U1/keyexpantion/SB0/n2799 ), .C(\U1/keyexpantion/SB0/n2579 ), .D(
        \U1/keyexpantion/SB0/n2578 ), .E(\U1/keyexpantion/SB0/n2577 ), .F(
        \U1/keyexpantion/SB0/n2576 ), .Y(\U1/keyexpantion/SB0/n2631 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U456  ( .A(\U1/keyexpantion/SB0/n2945 ), .B(\U1/keyexpantion/SB0/n2612 ), .Y(\U1/keyexpantion/SB0/n2747 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U455  ( .A(
        \U1/keyexpantion/SB0/n2874 ), .B(\U1/keyexpantion/SB0/n2962 ), .Y(
        \U1/keyexpantion/SB0/n2798 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U454  ( .A(
        \U1/keyexpantion/SB0/n2951 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2700 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U453  ( .A(\U1/keyexpantion/SB0/n2671 ), 
        .Y(\U1/keyexpantion/SB0/n2940 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U452  ( .A(
        \U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2723 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U451  ( .AN(
        \U1/keyexpantion/SB0/n2747 ), .B(\U1/keyexpantion/SB0/n2798 ), .C(
        \U1/keyexpantion/SB0/n2700 ), .D(\U1/keyexpantion/SB0/n2723 ), .Y(
        \U1/keyexpantion/SB0/n2586 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U450  ( .A(\U1/keyexpantion/SB0/n2932 ), .B(\U1/keyexpantion/SB0/n2782 ), .Y(\U1/keyexpantion/SB0/n2824 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U449  ( .A(
        \U1/keyexpantion/SB0/n2834 ), .B(\U1/keyexpantion/SB0/n2921 ), .Y(
        \U1/keyexpantion/SB0/n2680 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U448  ( .A0(
        \U1/keyexpantion/SB0/n2941 ), .A1(\U1/keyexpantion/SB0/n2840 ), .B0(
        \U1/keyexpantion/SB0/n2670 ), .Y(\U1/keyexpantion/SB0/n2580 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U447  ( .A(
        \U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2772 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U446  ( .AN(
        \U1/keyexpantion/SB0/n2824 ), .B(\U1/keyexpantion/SB0/n2680 ), .C(
        \U1/keyexpantion/SB0/n2580 ), .D(\U1/keyexpantion/SB0/n2772 ), .Y(
        \U1/keyexpantion/SB0/n2581 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U445  ( .A(\U1/keyexpantion/SB0/n2581 ), 
        .Y(\U1/keyexpantion/SB0/n2585 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U444  ( .A(\U1/keyexpantion/SB0/n2801 ), 
        .Y(\U1/keyexpantion/SB0/n2942 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U443  ( .A(\U1/keyexpantion/SB0/n2967 ), 
        .Y(\U1/keyexpantion/SB0/n2841 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U442  ( .A0(
        \U1/keyexpantion/SB0/n2962 ), .A1(\U1/keyexpantion/SB0/n2875 ), .B0(
        \U1/keyexpantion/SB0/n2942 ), .B1(\U1/keyexpantion/SB0/n2756 ), .C0(
        \U1/keyexpantion/SB0/n2841 ), .C1(\U1/keyexpantion/SB0/n2940 ), .Y(
        \U1/keyexpantion/SB0/n2584 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U441  ( .A0(
        \U1/keyexpantion/SB0/n2767 ), .A1(\U1/keyexpantion/SB0/n2945 ), .B0(
        \U1/keyexpantion/SB0/n2965 ), .B1(\U1/keyexpantion/SB0/n2966 ), .Y(
        \U1/keyexpantion/SB0/n2582 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U440  ( .A0(
        \U1/keyexpantion/SB0/n2818 ), .A1(\U1/keyexpantion/SB0/n2656 ), .B0(
        \U1/keyexpantion/SB0/n2874 ), .B1(\U1/keyexpantion/SB0/n2918 ), .C0(
        \U1/keyexpantion/SB0/n2582 ), .Y(\U1/keyexpantion/SB0/n2583 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U439  ( .AN(
        \U1/keyexpantion/SB0/n2586 ), .B(\U1/keyexpantion/SB0/n2585 ), .C(
        \U1/keyexpantion/SB0/n2584 ), .D(\U1/keyexpantion/SB0/n2583 ), .Y(
        \U1/keyexpantion/SB0/n2650 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U438  ( .A(\U1/keyexpantion/SB0/n2966 ), .B(\U1/keyexpantion/SB0/n2782 ), .Y(\U1/keyexpantion/SB0/n2665 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U437  ( .A0(
        \U1/keyexpantion/SB0/n2852 ), .A1(\U1/keyexpantion/SB0/n2966 ), .B0(
        \U1/keyexpantion/SB0/n2884 ), .Y(\U1/keyexpantion/SB0/n2591 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U436  ( .A(
        \U1/keyexpantion/SB0/n2884 ), .B(\U1/keyexpantion/SB0/n2872 ), .Y(
        \U1/keyexpantion/SB0/n2749 ) );
  AO22_X0P5M_A12TL \U1/keyexpantion/SB0/U435  ( .A0(
        \U1/keyexpantion/SB0/n2873 ), .A1(\U1/keyexpantion/SB0/n2656 ), .B0(
        \U1/keyexpantion/SB0/n2749 ), .B1(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2590 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U434  ( .A0(
        \U1/keyexpantion/SB0/n2927 ), .A1(\U1/keyexpantion/SB0/n2967 ), .B0(
        \U1/keyexpantion/SB0/n2671 ), .B1(\U1/keyexpantion/SB0/n2764 ), .C0(
        \U1/keyexpantion/SB0/n2929 ), .C1(\U1/keyexpantion/SB0/n2958 ), .Y(
        \U1/keyexpantion/SB0/n2589 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U433  ( .A(\U1/keyexpantion/SB0/n2767 ), 
        .Y(\U1/keyexpantion/SB0/n2835 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U432  ( .A(
        \U1/keyexpantion/SB0/n2960 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2861 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U431  ( .A(
        \U1/keyexpantion/SB0/n2834 ), .B(\U1/keyexpantion/SB0/n2656 ), .Y(
        \U1/keyexpantion/SB0/n2688 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U430  ( .A(
        \U1/keyexpantion/SB0/n2670 ), .B(\U1/keyexpantion/SB0/n2877 ), .Y(
        \U1/keyexpantion/SB0/n2708 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U429  ( .A(
        \U1/keyexpantion/SB0/n2834 ), .B(\U1/keyexpantion/SB0/n2875 ), .Y(
        \U1/keyexpantion/SB0/n2807 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U428  ( .A(
        \U1/keyexpantion/SB0/n2861 ), .B(\U1/keyexpantion/SB0/n2688 ), .C(
        \U1/keyexpantion/SB0/n2708 ), .D(\U1/keyexpantion/SB0/n2807 ), .Y(
        \U1/keyexpantion/SB0/n2588 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U427  ( .A(\U1/keyexpantion/SB0/n2854 ), .B(\U1/keyexpantion/SB0/n2767 ), .Y(\U1/keyexpantion/SB0/n2730 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U426  ( .A(
        \U1/keyexpantion/SB0/n2840 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2740 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U425  ( .A(
        \U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2756 ), .Y(
        \U1/keyexpantion/SB0/n2771 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U424  ( .AN(
        \U1/keyexpantion/SB0/n2730 ), .B(\U1/keyexpantion/SB0/n2740 ), .C(
        \U1/keyexpantion/SB0/n2771 ), .Y(\U1/keyexpantion/SB0/n2587 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U423  ( .A(\U1/keyexpantion/SB0/n2665 ), 
        .B(\U1/keyexpantion/SB0/n2591 ), .C(\U1/keyexpantion/SB0/n2590 ), .D(
        \U1/keyexpantion/SB0/n2589 ), .E(\U1/keyexpantion/SB0/n2588 ), .F(
        \U1/keyexpantion/SB0/n2587 ), .Y(\U1/keyexpantion/SB0/n2973 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U422  ( .A0(
        \U1/keyexpantion/SB0/n2670 ), .A1(\U1/keyexpantion/SB0/n2919 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2592 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U421  ( .A(
        \U1/keyexpantion/SB0/n2656 ), .B(\U1/keyexpantion/SB0/n2756 ), .Y(
        \U1/keyexpantion/SB0/n2793 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U420  ( .A(
        \U1/keyexpantion/SB0/n2873 ), .B(\U1/keyexpantion/SB0/n2942 ), .Y(
        \U1/keyexpantion/SB0/n2685 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U419  ( .A(
        \U1/keyexpantion/SB0/n2942 ), .B(\U1/keyexpantion/SB0/n2877 ), .Y(
        \U1/keyexpantion/SB0/n2736 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U418  ( .A(
        \U1/keyexpantion/SB0/n2592 ), .B(\U1/keyexpantion/SB0/n2793 ), .C(
        \U1/keyexpantion/SB0/n2685 ), .D(\U1/keyexpantion/SB0/n2736 ), .Y(
        \U1/keyexpantion/SB0/n2596 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U417  ( .A0(
        \U1/keyexpantion/SB0/n2945 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2671 ), .B1(\U1/keyexpantion/SB0/n2917 ), .C0(
        \U1/keyexpantion/SB0/n2946 ), .C1(\U1/keyexpantion/SB0/n2782 ), .Y(
        \U1/keyexpantion/SB0/n2595 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U416  ( .A(
        \U1/keyexpantion/SB0/n2876 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2717 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U415  ( .A(
        \U1/keyexpantion/SB0/n2875 ), .B(\U1/keyexpantion/SB0/n2948 ), .Y(
        \U1/keyexpantion/SB0/n2857 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U414  ( .A(
        \U1/keyexpantion/SB0/n2875 ), .B(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2704 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U413  ( .A(
        \U1/keyexpantion/SB0/n2951 ), .B(\U1/keyexpantion/SB0/n2941 ), .Y(
        \U1/keyexpantion/SB0/n2666 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U412  ( .A(
        \U1/keyexpantion/SB0/n2717 ), .B(\U1/keyexpantion/SB0/n2857 ), .C(
        \U1/keyexpantion/SB0/n2704 ), .D(\U1/keyexpantion/SB0/n2666 ), .Y(
        \U1/keyexpantion/SB0/n2594 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U411  ( .A(
        \U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2779 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U410  ( .A(
        \U1/keyexpantion/SB0/n2960 ), .B(\U1/keyexpantion/SB0/n2921 ), .Y(
        \U1/keyexpantion/SB0/n2752 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U409  ( .A(
        \U1/keyexpantion/SB0/n2950 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2803 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U408  ( .A(
        \U1/keyexpantion/SB0/n2682 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2653 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U407  ( .A(
        \U1/keyexpantion/SB0/n2779 ), .B(\U1/keyexpantion/SB0/n2752 ), .C(
        \U1/keyexpantion/SB0/n2803 ), .D(\U1/keyexpantion/SB0/n2653 ), .Y(
        \U1/keyexpantion/SB0/n2593 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U406  ( .A(\U1/keyexpantion/SB0/n2596 ), 
        .B(\U1/keyexpantion/SB0/n2595 ), .C(\U1/keyexpantion/SB0/n2594 ), .D(
        \U1/keyexpantion/SB0/n2593 ), .Y(\U1/keyexpantion/SB0/n2639 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U405  ( .A(\U1/keyexpantion/SB0/n2631 ), 
        .B(\U1/keyexpantion/SB0/n2650 ), .C(\U1/keyexpantion/SB0/n2973 ), .D(
        \U1/keyexpantion/SB0/n2639 ), .Y(\U1/keyexpantion/SB0/n2606 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U404  ( .A(\U1/keyexpantion/SB0/n2927 ), 
        .Y(\U1/keyexpantion/SB0/n2830 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U403  ( .A0(
        \U1/keyexpantion/SB0/n2782 ), .A1(\U1/keyexpantion/SB0/n2613 ), .B0(
        \U1/keyexpantion/SB0/n2751 ), .B1(\U1/keyexpantion/SB0/n2958 ), .Y(
        \U1/keyexpantion/SB0/n2597 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U402  ( .A0(
        \U1/keyexpantion/SB0/n2830 ), .A1(\U1/keyexpantion/SB0/n2882 ), .B0(
        \U1/keyexpantion/SB0/n2952 ), .B1(\U1/keyexpantion/SB0/n2960 ), .C0(
        \U1/keyexpantion/SB0/n2597 ), .Y(\U1/keyexpantion/SB0/n2605 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U401  ( .A(
        \U1/keyexpantion/SB0/n2851 ), .B(\U1/keyexpantion/SB0/n2854 ), .Y(
        \U1/keyexpantion/SB0/n2850 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U400  ( .A0(
        \U1/keyexpantion/SB0/n2785 ), .A1(\U1/keyexpantion/SB0/n2854 ), .B0(
        \U1/keyexpantion/SB0/n2767 ), .B1(\U1/keyexpantion/SB0/n2916 ), .Y(
        \U1/keyexpantion/SB0/n2598 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U399  ( .A0(
        \U1/keyexpantion/SB0/n2682 ), .A1(\U1/keyexpantion/SB0/n2850 ), .B0(
        \U1/keyexpantion/SB0/n2922 ), .B1(\U1/keyexpantion/SB0/n2941 ), .C0(
        \U1/keyexpantion/SB0/n2598 ), .Y(\U1/keyexpantion/SB0/n2604 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U398  ( .A(
        \U1/keyexpantion/SB0/n2946 ), .B(\U1/keyexpantion/SB0/n2784 ), .Y(
        \U1/keyexpantion/SB0/n2602 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U397  ( .A(\U1/keyexpantion/SB0/n2875 ), .B(\U1/keyexpantion/SB0/n2921 ), .Y(\U1/keyexpantion/SB0/n2842 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U396  ( .A(\U1/keyexpantion/SB0/n2842 ), 
        .Y(\U1/keyexpantion/SB0/n2601 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U395  ( .A(\U1/keyexpantion/SB0/n2833 ), .B(\U1/keyexpantion/SB0/n2927 ), .Y(\U1/keyexpantion/SB0/n2714 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U394  ( .A(\U1/keyexpantion/SB0/n2932 ), .B(\U1/keyexpantion/SB0/n2930 ), .Y(\U1/keyexpantion/SB0/n2867 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U393  ( .A(\U1/keyexpantion/SB0/n2867 ), 
        .Y(\U1/keyexpantion/SB0/n2599 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U392  ( .A(
        \U1/keyexpantion/SB0/n2882 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2724 ) );
  NAND3B_X0P5M_A12TL \U1/keyexpantion/SB0/U391  ( .AN(
        \U1/keyexpantion/SB0/n2714 ), .B(\U1/keyexpantion/SB0/n2599 ), .C(
        \U1/keyexpantion/SB0/n2724 ), .Y(\U1/keyexpantion/SB0/n2600 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U390  ( .A0(
        \U1/keyexpantion/SB0/n2841 ), .A1(\U1/keyexpantion/SB0/n2602 ), .B0(
        \U1/keyexpantion/SB0/n2818 ), .B1(\U1/keyexpantion/SB0/n2601 ), .C0(
        \U1/keyexpantion/SB0/n2600 ), .Y(\U1/keyexpantion/SB0/n2603 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U389  ( .AN(
        \U1/keyexpantion/SB0/n2606 ), .B(\U1/keyexpantion/SB0/n2605 ), .C(
        \U1/keyexpantion/SB0/n2604 ), .D(\U1/keyexpantion/SB0/n2603 ), .Y(
        \U1/keyexpantion/ws [24]) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U388  ( .A(\U1/keyexpantion/SB0/n2854 ), .B(\U1/keyexpantion/SB0/n2671 ), .Y(\U1/keyexpantion/SB0/n2731 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U387  ( .A(\U1/keyexpantion/SB0/n2801 ), .B(\U1/keyexpantion/SB0/n2851 ), .Y(\U1/keyexpantion/SB0/n2691 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U386  ( .A(\U1/keyexpantion/SB0/n2818 ), .B(\U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2800 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U385  ( .A0(
        \U1/keyexpantion/SB0/n2800 ), .A1(\U1/keyexpantion/SB0/n2854 ), .B0(
        \U1/keyexpantion/SB0/n2964 ), .Y(\U1/keyexpantion/SB0/n2611 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U384  ( .A(
        \U1/keyexpantion/SB0/n2882 ), .B(\U1/keyexpantion/SB0/n2951 ), .Y(
        \U1/keyexpantion/SB0/n2707 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U383  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2882 ), .Y(
        \U1/keyexpantion/SB0/n2806 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U382  ( .A(
        \U1/keyexpantion/SB0/n2948 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2739 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U381  ( .A(
        \U1/keyexpantion/SB0/n2707 ), .B(\U1/keyexpantion/SB0/n2806 ), .C(
        \U1/keyexpantion/SB0/n2739 ), .Y(\U1/keyexpantion/SB0/n2610 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U380  ( .A(\U1/keyexpantion/SB0/n2882 ), .B(\U1/keyexpantion/SB0/n2962 ), .Y(\U1/keyexpantion/SB0/n2766 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U379  ( .A(\U1/keyexpantion/SB0/n2948 ), .B(\U1/keyexpantion/SB0/n2939 ), .C(\U1/keyexpantion/SB0/n2960 ), .Y(
        \U1/keyexpantion/SB0/n2607 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U378  ( .A0(
        \U1/keyexpantion/SB0/n2766 ), .A1(\U1/keyexpantion/SB0/n2928 ), .B0(
        \U1/keyexpantion/SB0/n2607 ), .B1(\U1/keyexpantion/SB0/n2958 ), .C0(
        \U1/keyexpantion/SB0/n2801 ), .C1(\U1/keyexpantion/SB0/n2833 ), .Y(
        \U1/keyexpantion/SB0/n2609 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U377  ( .A0(
        \U1/keyexpantion/SB0/n2929 ), .A1(\U1/keyexpantion/SB0/n2957 ), .B0(
        \U1/keyexpantion/SB0/n2930 ), .B1(\U1/keyexpantion/SB0/n2927 ), .Y(
        \U1/keyexpantion/SB0/n2608 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U376  ( .A(\U1/keyexpantion/SB0/n2731 ), 
        .B(\U1/keyexpantion/SB0/n2691 ), .C(\U1/keyexpantion/SB0/n2611 ), .D(
        \U1/keyexpantion/SB0/n2610 ), .E(\U1/keyexpantion/SB0/n2609 ), .F(
        \U1/keyexpantion/SB0/n2608 ), .Y(\U1/keyexpantion/SB0/n2972 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U375  ( .A(\U1/keyexpantion/SB0/n2782 ), .B(\U1/keyexpantion/SB0/n2767 ), .Y(\U1/keyexpantion/SB0/n2657 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U374  ( .A0(
        \U1/keyexpantion/SB0/n2782 ), .A1(\U1/keyexpantion/SB0/n2872 ), .B0(
        \U1/keyexpantion/SB0/n2671 ), .Y(\U1/keyexpantion/SB0/n2618 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U373  ( .A(\U1/keyexpantion/SB0/n2876 ), .B(\U1/keyexpantion/SB0/n2882 ), .Y(\U1/keyexpantion/SB0/n2659 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U372  ( .A0(
        \U1/keyexpantion/SB0/n2764 ), .A1(\U1/keyexpantion/SB0/n2932 ), .B0(
        \U1/keyexpantion/SB0/n2659 ), .B1(\U1/keyexpantion/SB0/n2946 ), .Y(
        \U1/keyexpantion/SB0/n2617 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U371  ( .A0(
        \U1/keyexpantion/SB0/n2751 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2916 ), .B1(\U1/keyexpantion/SB0/n2801 ), .C0(
        \U1/keyexpantion/SB0/n2930 ), .C1(\U1/keyexpantion/SB0/n2852 ), .Y(
        \U1/keyexpantion/SB0/n2616 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U370  ( .A(\U1/keyexpantion/SB0/n2965 ), .B(\U1/keyexpantion/SB0/n2612 ), .Y(\U1/keyexpantion/SB0/n2715 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U369  ( .A(
        \U1/keyexpantion/SB0/n2952 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2722 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U368  ( .A(
        \U1/keyexpantion/SB0/n2873 ), .B(\U1/keyexpantion/SB0/n2947 ), .Y(
        \U1/keyexpantion/SB0/n2732 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U367  ( .A(
        \U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2962 ), .Y(
        \U1/keyexpantion/SB0/n2836 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U366  ( .AN(
        \U1/keyexpantion/SB0/n2715 ), .B(\U1/keyexpantion/SB0/n2722 ), .C(
        \U1/keyexpantion/SB0/n2732 ), .D(\U1/keyexpantion/SB0/n2836 ), .Y(
        \U1/keyexpantion/SB0/n2615 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U365  ( .A(\U1/keyexpantion/SB0/n2833 ), .B(\U1/keyexpantion/SB0/n2613 ), .Y(\U1/keyexpantion/SB0/n2815 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U364  ( .A(\U1/keyexpantion/SB0/n2932 ), .B(\U1/keyexpantion/SB0/n2916 ), .Y(\U1/keyexpantion/SB0/n2868 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U362  ( .A(
        \U1/keyexpantion/SB0/n2656 ), .B(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2681 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U360  ( .A(\U1/keyexpantion/SB0/n2657 ), 
        .B(\U1/keyexpantion/SB0/n2618 ), .C(\U1/keyexpantion/SB0/n2617 ), .D(
        \U1/keyexpantion/SB0/n2616 ), .E(\U1/keyexpantion/SB0/n2615 ), .F(
        \U1/keyexpantion/SB0/n2614 ), .Y(\U1/keyexpantion/SB0/n2651 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U359  ( .A(\U1/keyexpantion/SB0/n2849 ), .B(\U1/keyexpantion/SB0/n2671 ), .Y(\U1/keyexpantion/SB0/n2669 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U358  ( .A(\U1/keyexpantion/SB0/n2801 ), .B(\U1/keyexpantion/SB0/n2751 ), .Y(\U1/keyexpantion/SB0/n2881 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U357  ( .A(\U1/keyexpantion/SB0/n2782 ), .B(\U1/keyexpantion/SB0/n2852 ), .Y(\U1/keyexpantion/SB0/n2719 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U356  ( .A(\U1/keyexpantion/SB0/n2967 ), .B(\U1/keyexpantion/SB0/n2852 ), .Y(\U1/keyexpantion/SB0/n2734 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U355  ( .A(
        \U1/keyexpantion/SB0/n2877 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2794 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U354  ( .A(
        \U1/keyexpantion/SB0/n2948 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2686 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U353  ( .A(
        \U1/keyexpantion/SB0/n2952 ), .B(\U1/keyexpantion/SB0/n2948 ), .Y(
        \U1/keyexpantion/SB0/n2780 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U352  ( .A(
        \U1/keyexpantion/SB0/n2841 ), .B(\U1/keyexpantion/SB0/n2919 ), .Y(
        \U1/keyexpantion/SB0/n2705 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U351  ( .A(
        \U1/keyexpantion/SB0/n2794 ), .B(\U1/keyexpantion/SB0/n2686 ), .C(
        \U1/keyexpantion/SB0/n2780 ), .D(\U1/keyexpantion/SB0/n2705 ), .Y(
        \U1/keyexpantion/SB0/n2622 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U350  ( .A(\U1/keyexpantion/SB0/n2967 ), .B(\U1/keyexpantion/SB0/n2767 ), .Y(\U1/keyexpantion/SB0/n2755 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U349  ( .A(\U1/keyexpantion/SB0/n2966 ), .B(\U1/keyexpantion/SB0/n2751 ), .Y(\U1/keyexpantion/SB0/n2855 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U348  ( .A(\U1/keyexpantion/SB0/n2872 ), .B(\U1/keyexpantion/SB0/n2932 ), .Y(\U1/keyexpantion/SB0/n2805 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U347  ( .A(\U1/keyexpantion/SB0/n2833 ), .B(\U1/keyexpantion/SB0/n2932 ), .Y(\U1/keyexpantion/SB0/n2655 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U346  ( .A0(
        \U1/keyexpantion/SB0/n2932 ), .A1(\U1/keyexpantion/SB0/n2967 ), .B0(
        \U1/keyexpantion/SB0/n2767 ), .B1(\U1/keyexpantion/SB0/n2872 ), .Y(
        \U1/keyexpantion/SB0/n2620 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U345  ( .A0(
        \U1/keyexpantion/SB0/n2751 ), .A1(\U1/keyexpantion/SB0/n2964 ), .B0(
        \U1/keyexpantion/SB0/n2764 ), .B1(\U1/keyexpantion/SB0/n2801 ), .Y(
        \U1/keyexpantion/SB0/n2619 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U344  ( .A(\U1/keyexpantion/SB0/n2755 ), 
        .B(\U1/keyexpantion/SB0/n2855 ), .C(\U1/keyexpantion/SB0/n2805 ), .D(
        \U1/keyexpantion/SB0/n2655 ), .E(\U1/keyexpantion/SB0/n2620 ), .F(
        \U1/keyexpantion/SB0/n2619 ), .Y(\U1/keyexpantion/SB0/n2621 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U343  ( .A(\U1/keyexpantion/SB0/n2669 ), 
        .B(\U1/keyexpantion/SB0/n2881 ), .C(\U1/keyexpantion/SB0/n2719 ), .D(
        \U1/keyexpantion/SB0/n2734 ), .E(\U1/keyexpantion/SB0/n2622 ), .F(
        \U1/keyexpantion/SB0/n2621 ), .Y(\U1/keyexpantion/SB0/n2640 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U342  ( .A0(
        \U1/keyexpantion/SB0/n2877 ), .A1(\U1/keyexpantion/SB0/n2874 ), .B0(
        \U1/keyexpantion/SB0/n2951 ), .B1(\U1/keyexpantion/SB0/n2818 ), .C0(
        \U1/keyexpantion/SB0/n2640 ), .Y(\U1/keyexpantion/SB0/n2623 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U341  ( .A(\U1/keyexpantion/SB0/n2623 ), 
        .Y(\U1/keyexpantion/SB0/n2630 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U340  ( .A(
        \U1/keyexpantion/SB0/n2930 ), .B(\U1/keyexpantion/SB0/n2872 ), .Y(
        \U1/keyexpantion/SB0/n2920 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U339  ( .A0(
        \U1/keyexpantion/SB0/n2876 ), .A1(\U1/keyexpantion/SB0/n2920 ), .B0(
        \U1/keyexpantion/SB0/n2952 ), .Y(\U1/keyexpantion/SB0/n2626 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U338  ( .A0(
        \U1/keyexpantion/SB0/n2841 ), .A1(\U1/keyexpantion/SB0/n2941 ), .B0(
        \U1/keyexpantion/SB0/n2883 ), .Y(\U1/keyexpantion/SB0/n2625 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U337  ( .A0(
        \U1/keyexpantion/SB0/n2840 ), .A1(\U1/keyexpantion/SB0/n2882 ), .B0(
        \U1/keyexpantion/SB0/n2947 ), .Y(\U1/keyexpantion/SB0/n2624 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U336  ( .A(
        \U1/keyexpantion/SB0/n2873 ), .B(\U1/keyexpantion/SB0/n2940 ), .Y(
        \U1/keyexpantion/SB0/n2698 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U335  ( .A(
        \U1/keyexpantion/SB0/n2626 ), .B(\U1/keyexpantion/SB0/n2625 ), .C(
        \U1/keyexpantion/SB0/n2624 ), .D(\U1/keyexpantion/SB0/n2698 ), .Y(
        \U1/keyexpantion/SB0/n2629 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U334  ( .A(\U1/keyexpantion/SB0/n2939 ), .B(\U1/keyexpantion/SB0/n2834 ), .Y(\U1/keyexpantion/SB0/n2888 ) );
  AND3_X0P5M_A12TL \U1/keyexpantion/SB0/U333  ( .A(\U1/keyexpantion/SB0/n2888 ), .B(\U1/keyexpantion/SB0/n2929 ), .C(\U1/keyexpantion/SB0/n2916 ), .Y(
        \U1/keyexpantion/SB0/n2627 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U332  ( .A0(
        \U1/keyexpantion/SB0/n2872 ), .A1(\U1/keyexpantion/SB0/n2966 ), .B0(
        \U1/keyexpantion/SB0/n2627 ), .B1(\U1/keyexpantion/SB0/n2927 ), .C0(
        \U1/keyexpantion/SB0/n2965 ), .C1(\U1/keyexpantion/SB0/n2957 ), .Y(
        \U1/keyexpantion/SB0/n2628 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U331  ( .A(\U1/keyexpantion/SB0/n2972 ), 
        .B(\U1/keyexpantion/SB0/n2651 ), .C(\U1/keyexpantion/SB0/n2631 ), .D(
        \U1/keyexpantion/SB0/n2630 ), .E(\U1/keyexpantion/SB0/n2629 ), .F(
        \U1/keyexpantion/SB0/n2628 ), .Y(\U1/keyexpantion/ws [25]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U330  ( .A0(
        \U1/keyexpantion/SB0/n2921 ), .A1(\U1/keyexpantion/SB0/n2941 ), .B0(
        \U1/keyexpantion/SB0/n2962 ), .B1(\U1/keyexpantion/SB0/n2952 ), .Y(
        \U1/keyexpantion/SB0/n2632 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U329  ( .A0(
        \U1/keyexpantion/SB0/n2851 ), .A1(\U1/keyexpantion/SB0/n2966 ), .B0(
        \U1/keyexpantion/SB0/n2801 ), .B1(\U1/keyexpantion/SB0/n2872 ), .C0(
        \U1/keyexpantion/SB0/n2632 ), .Y(\U1/keyexpantion/SB0/n2638 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U328  ( .A(
        \U1/keyexpantion/SB0/n2947 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2735 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U327  ( .A(
        \U1/keyexpantion/SB0/n2921 ), .B(\U1/keyexpantion/SB0/n2876 ), .Y(
        \U1/keyexpantion/SB0/n2716 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U326  ( .A(
        \U1/keyexpantion/SB0/n2941 ), .B(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2684 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U325  ( .A(
        \U1/keyexpantion/SB0/n2840 ), .B(\U1/keyexpantion/SB0/n2883 ), .Y(
        \U1/keyexpantion/SB0/n2703 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U324  ( .A(
        \U1/keyexpantion/SB0/n2735 ), .B(\U1/keyexpantion/SB0/n2716 ), .C(
        \U1/keyexpantion/SB0/n2684 ), .D(\U1/keyexpantion/SB0/n2703 ), .Y(
        \U1/keyexpantion/SB0/n2637 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U323  ( .A(
        \U1/keyexpantion/SB0/n2967 ), .B(\U1/keyexpantion/SB0/n2945 ), .Y(
        \U1/keyexpantion/SB0/n2829 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U322  ( .A0(
        \U1/keyexpantion/SB0/n2877 ), .A1(\U1/keyexpantion/SB0/n2829 ), .B0(
        \U1/keyexpantion/SB0/n2951 ), .Y(\U1/keyexpantion/SB0/n2635 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U321  ( .A0(
        \U1/keyexpantion/SB0/n2948 ), .A1(\U1/keyexpantion/SB0/n2818 ), .B0(
        \U1/keyexpantion/SB0/n2830 ), .Y(\U1/keyexpantion/SB0/n2634 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U320  ( .A0(
        \U1/keyexpantion/SB0/n2835 ), .A1(\U1/keyexpantion/SB0/n2875 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2633 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U319  ( .A(
        \U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2948 ), .Y(
        \U1/keyexpantion/SB0/n2802 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U318  ( .A(
        \U1/keyexpantion/SB0/n2635 ), .B(\U1/keyexpantion/SB0/n2634 ), .C(
        \U1/keyexpantion/SB0/n2633 ), .D(\U1/keyexpantion/SB0/n2802 ), .Y(
        \U1/keyexpantion/SB0/n2636 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U317  ( .A(\U1/keyexpantion/SB0/n2641 ), 
        .B(\U1/keyexpantion/SB0/n2640 ), .C(\U1/keyexpantion/SB0/n2639 ), .D(
        \U1/keyexpantion/SB0/n2638 ), .E(\U1/keyexpantion/SB0/n2637 ), .F(
        \U1/keyexpantion/SB0/n2636 ), .Y(\U1/keyexpantion/SB0/n2971 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U316  ( .A0(
        \U1/keyexpantion/SB0/n2756 ), .A1(\U1/keyexpantion/SB0/n2952 ), .B0(
        \U1/keyexpantion/SB0/n2960 ), .B1(\U1/keyexpantion/SB0/n2874 ), .C0(
        \U1/keyexpantion/SB0/n2971 ), .Y(\U1/keyexpantion/SB0/n2642 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U315  ( .A(\U1/keyexpantion/SB0/n2642 ), 
        .Y(\U1/keyexpantion/SB0/n2649 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U314  ( .A(\U1/keyexpantion/SB0/n2883 ), .B(\U1/keyexpantion/SB0/n2670 ), .Y(\U1/keyexpantion/SB0/n2792 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U313  ( .A1N(
        \U1/keyexpantion/SB0/n2792 ), .A0(\U1/keyexpantion/SB0/n2922 ), .B0(
        \U1/keyexpantion/SB0/n2873 ), .Y(\U1/keyexpantion/SB0/n2645 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U312  ( .A0(
        \U1/keyexpantion/SB0/n2841 ), .A1(\U1/keyexpantion/SB0/n2749 ), .B0(
        \U1/keyexpantion/SB0/n2921 ), .Y(\U1/keyexpantion/SB0/n2644 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U311  ( .A0(
        \U1/keyexpantion/SB0/n2948 ), .A1(\U1/keyexpantion/SB0/n2882 ), .B0(
        \U1/keyexpantion/SB0/n2942 ), .Y(\U1/keyexpantion/SB0/n2643 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U310  ( .A(
        \U1/keyexpantion/SB0/n2919 ), .B(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2699 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U309  ( .A(
        \U1/keyexpantion/SB0/n2645 ), .B(\U1/keyexpantion/SB0/n2644 ), .C(
        \U1/keyexpantion/SB0/n2643 ), .D(\U1/keyexpantion/SB0/n2699 ), .Y(
        \U1/keyexpantion/SB0/n2648 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U308  ( .A(\U1/keyexpantion/SB0/n2918 ), .B(\U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2949 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U307  ( .A(\U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2875 ), .Y(\U1/keyexpantion/SB0/n2646 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U306  ( .A0(
        \U1/keyexpantion/SB0/n2949 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2646 ), .B1(\U1/keyexpantion/SB0/n2930 ), .C0(
        \U1/keyexpantion/SB0/n2852 ), .C1(\U1/keyexpantion/SB0/n2854 ), .Y(
        \U1/keyexpantion/SB0/n2647 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U305  ( .A(\U1/keyexpantion/SB0/n2652 ), 
        .B(\U1/keyexpantion/SB0/n2651 ), .C(\U1/keyexpantion/SB0/n2650 ), .D(
        \U1/keyexpantion/SB0/n2649 ), .E(\U1/keyexpantion/SB0/n2648 ), .F(
        \U1/keyexpantion/SB0/n2647 ), .Y(\U1/keyexpantion/ws [26]) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U304  ( .A(
        \U1/keyexpantion/SB0/n2756 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2954 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U303  ( .AN(
        \U1/keyexpantion/SB0/n2655 ), .B(\U1/keyexpantion/SB0/n2654 ), .C(
        \U1/keyexpantion/SB0/n2653 ), .D(\U1/keyexpantion/SB0/n2954 ), .Y(
        \U1/keyexpantion/SB0/n2662 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U302  ( .A0(
        \U1/keyexpantion/SB0/n2656 ), .A1(\U1/keyexpantion/SB0/n2921 ), .B0(
        \U1/keyexpantion/SB0/n2818 ), .Y(\U1/keyexpantion/SB0/n2658 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U299  ( .A(\U1/keyexpantion/SB0/n2874 ), .B(\U1/keyexpantion/SB0/n2942 ), .Y(\U1/keyexpantion/SB0/n2885 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U298  ( .A0(
        \U1/keyexpantion/SB0/n2764 ), .A1(\U1/keyexpantion/SB0/n2964 ), .B0(
        \U1/keyexpantion/SB0/n2885 ), .B1(\U1/keyexpantion/SB0/n2917 ), .C0(
        \U1/keyexpantion/SB0/n2958 ), .C1(\U1/keyexpantion/SB0/n2967 ), .Y(
        \U1/keyexpantion/SB0/n2660 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U297  ( .A(\U1/keyexpantion/SB0/n2665 ), 
        .B(\U1/keyexpantion/SB0/n2664 ), .C(\U1/keyexpantion/SB0/n2663 ), .D(
        \U1/keyexpantion/SB0/n2662 ), .E(\U1/keyexpantion/SB0/n2661 ), .F(
        \U1/keyexpantion/SB0/n2660 ), .Y(\U1/keyexpantion/SB0/n2848 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U296  ( .AN(
        \U1/keyexpantion/SB0/n2669 ), .B(\U1/keyexpantion/SB0/n2668 ), .C(
        \U1/keyexpantion/SB0/n2667 ), .D(\U1/keyexpantion/SB0/n2666 ), .Y(
        \U1/keyexpantion/SB0/n2679 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U295  ( .A0(
        \U1/keyexpantion/SB0/n2952 ), .A1(\U1/keyexpantion/SB0/n2841 ), .B0(
        \U1/keyexpantion/SB0/n2947 ), .B1(\U1/keyexpantion/SB0/n2840 ), .C0(
        \U1/keyexpantion/SB0/n2670 ), .C1(\U1/keyexpantion/SB0/n2962 ), .Y(
        \U1/keyexpantion/SB0/n2678 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U294  ( .A0(
        \U1/keyexpantion/SB0/n2916 ), .A1(\U1/keyexpantion/SB0/n2801 ), .B0(
        \U1/keyexpantion/SB0/n2671 ), .B1(\U1/keyexpantion/SB0/n2764 ), .Y(
        \U1/keyexpantion/SB0/n2672 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U293  ( .A0(
        \U1/keyexpantion/SB0/n2818 ), .A1(\U1/keyexpantion/SB0/n2835 ), .B0(
        \U1/keyexpantion/SB0/n2834 ), .B1(\U1/keyexpantion/SB0/n2919 ), .C0(
        \U1/keyexpantion/SB0/n2672 ), .Y(\U1/keyexpantion/SB0/n2677 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U292  ( .A(
        \U1/keyexpantion/SB0/n2927 ), .B(\U1/keyexpantion/SB0/n2966 ), .Y(
        \U1/keyexpantion/SB0/n2674 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U291  ( .A0(
        \U1/keyexpantion/SB0/n2756 ), .A1(\U1/keyexpantion/SB0/n2675 ), .B0(
        \U1/keyexpantion/SB0/n2948 ), .B1(\U1/keyexpantion/SB0/n2674 ), .C0(
        \U1/keyexpantion/SB0/n2673 ), .Y(\U1/keyexpantion/SB0/n2676 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U290  ( .AN(
        \U1/keyexpantion/SB0/n2679 ), .B(\U1/keyexpantion/SB0/n2678 ), .C(
        \U1/keyexpantion/SB0/n2677 ), .D(\U1/keyexpantion/SB0/n2676 ), .Y(
        \U1/keyexpantion/SB0/n2893 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U289  ( .A(\U1/keyexpantion/SB0/n2680 ), 
        .Y(\U1/keyexpantion/SB0/n2696 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U288  ( .A0(
        \U1/keyexpantion/SB0/n2785 ), .A1(\U1/keyexpantion/SB0/n2854 ), .B0(
        \U1/keyexpantion/SB0/n2681 ), .Y(\U1/keyexpantion/SB0/n2695 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U287  ( .A0(
        \U1/keyexpantion/SB0/n2948 ), .A1(\U1/keyexpantion/SB0/n2947 ), .B0(
        \U1/keyexpantion/SB0/n2918 ), .B1(\U1/keyexpantion/SB0/n2682 ), .Y(
        \U1/keyexpantion/SB0/n2683 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U286  ( .A0(
        \U1/keyexpantion/SB0/n2929 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2945 ), .B1(\U1/keyexpantion/SB0/n2957 ), .C0(
        \U1/keyexpantion/SB0/n2683 ), .Y(\U1/keyexpantion/SB0/n2694 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U285  ( .A(
        \U1/keyexpantion/SB0/n2687 ), .B(\U1/keyexpantion/SB0/n2686 ), .C(
        \U1/keyexpantion/SB0/n2685 ), .D(\U1/keyexpantion/SB0/n2684 ), .Y(
        \U1/keyexpantion/SB0/n2693 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U284  ( .AN(
        \U1/keyexpantion/SB0/n2691 ), .B(\U1/keyexpantion/SB0/n2690 ), .C(
        \U1/keyexpantion/SB0/n2689 ), .D(\U1/keyexpantion/SB0/n2688 ), .Y(
        \U1/keyexpantion/SB0/n2692 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U283  ( .A(\U1/keyexpantion/SB0/n2697 ), 
        .B(\U1/keyexpantion/SB0/n2696 ), .C(\U1/keyexpantion/SB0/n2695 ), .D(
        \U1/keyexpantion/SB0/n2694 ), .E(\U1/keyexpantion/SB0/n2693 ), .F(
        \U1/keyexpantion/SB0/n2692 ), .Y(\U1/keyexpantion/SB0/n2797 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U282  ( .A0(
        \U1/keyexpantion/SB0/n2884 ), .A1(\U1/keyexpantion/SB0/n2801 ), .B0(
        \U1/keyexpantion/SB0/n2698 ), .Y(\U1/keyexpantion/SB0/n2713 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U281  ( .AN(
        \U1/keyexpantion/SB0/n2702 ), .B(\U1/keyexpantion/SB0/n2701 ), .C(
        \U1/keyexpantion/SB0/n2700 ), .D(\U1/keyexpantion/SB0/n2699 ), .Y(
        \U1/keyexpantion/SB0/n2712 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U280  ( .A(
        \U1/keyexpantion/SB0/n2939 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2953 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U279  ( .A(
        \U1/keyexpantion/SB0/n2705 ), .B(\U1/keyexpantion/SB0/n2704 ), .C(
        \U1/keyexpantion/SB0/n2703 ), .D(\U1/keyexpantion/SB0/n2953 ), .Y(
        \U1/keyexpantion/SB0/n2711 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U278  ( .A(
        \U1/keyexpantion/SB0/n2709 ), .B(\U1/keyexpantion/SB0/n2708 ), .C(
        \U1/keyexpantion/SB0/n2707 ), .D(\U1/keyexpantion/SB0/n2706 ), .Y(
        \U1/keyexpantion/SB0/n2710 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U277  ( .A(\U1/keyexpantion/SB0/n2715 ), 
        .B(\U1/keyexpantion/SB0/n2714 ), .C(\U1/keyexpantion/SB0/n2713 ), .D(
        \U1/keyexpantion/SB0/n2712 ), .E(\U1/keyexpantion/SB0/n2711 ), .F(
        \U1/keyexpantion/SB0/n2710 ), .Y(\U1/keyexpantion/SB0/n2821 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U276  ( .AN(
        \U1/keyexpantion/SB0/n2719 ), .B(\U1/keyexpantion/SB0/n2718 ), .C(
        \U1/keyexpantion/SB0/n2717 ), .D(\U1/keyexpantion/SB0/n2716 ), .Y(
        \U1/keyexpantion/SB0/n2728 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U275  ( .A(
        \U1/keyexpantion/SB0/n2723 ), .B(\U1/keyexpantion/SB0/n2722 ), .C(
        \U1/keyexpantion/SB0/n2721 ), .D(\U1/keyexpantion/SB0/n2720 ), .Y(
        \U1/keyexpantion/SB0/n2727 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U274  ( .A(\U1/keyexpantion/SB0/n2883 ), .B(\U1/keyexpantion/SB0/n2940 ), .C(\U1/keyexpantion/SB0/n2942 ), .Y(
        \U1/keyexpantion/SB0/n2725 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U273  ( .A0(
        \U1/keyexpantion/SB0/n2725 ), .A1(\U1/keyexpantion/SB0/n2930 ), .B0(
        \U1/keyexpantion/SB0/n2764 ), .B1(\U1/keyexpantion/SB0/n2966 ), .C0(
        \U1/keyexpantion/SB0/n2724 ), .Y(\U1/keyexpantion/SB0/n2726 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U272  ( .A(\U1/keyexpantion/SB0/n2731 ), 
        .B(\U1/keyexpantion/SB0/n2730 ), .C(\U1/keyexpantion/SB0/n2729 ), .D(
        \U1/keyexpantion/SB0/n2728 ), .E(\U1/keyexpantion/SB0/n2727 ), .F(
        \U1/keyexpantion/SB0/n2726 ), .Y(\U1/keyexpantion/SB0/n2869 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U271  ( .A0(
        \U1/keyexpantion/SB0/n2764 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2732 ), .Y(\U1/keyexpantion/SB0/n2746 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U270  ( .A0(
        \U1/keyexpantion/SB0/n2873 ), .A1(\U1/keyexpantion/SB0/n2875 ), .B0(
        \U1/keyexpantion/SB0/n2951 ), .B1(\U1/keyexpantion/SB0/n2840 ), .Y(
        \U1/keyexpantion/SB0/n2733 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U269  ( .A0(
        \U1/keyexpantion/SB0/n2784 ), .A1(\U1/keyexpantion/SB0/n2872 ), .B0(
        \U1/keyexpantion/SB0/n2785 ), .B1(\U1/keyexpantion/SB0/n2849 ), .C0(
        \U1/keyexpantion/SB0/n2733 ), .Y(\U1/keyexpantion/SB0/n2745 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U268  ( .A(\U1/keyexpantion/SB0/n2734 ), 
        .Y(\U1/keyexpantion/SB0/n2737 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U267  ( .AN(
        \U1/keyexpantion/SB0/n2738 ), .B(\U1/keyexpantion/SB0/n2737 ), .C(
        \U1/keyexpantion/SB0/n2736 ), .D(\U1/keyexpantion/SB0/n2735 ), .Y(
        \U1/keyexpantion/SB0/n2744 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U266  ( .A(
        \U1/keyexpantion/SB0/n2742 ), .B(\U1/keyexpantion/SB0/n2741 ), .C(
        \U1/keyexpantion/SB0/n2740 ), .D(\U1/keyexpantion/SB0/n2739 ), .Y(
        \U1/keyexpantion/SB0/n2743 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U265  ( .A(\U1/keyexpantion/SB0/n2748 ), 
        .B(\U1/keyexpantion/SB0/n2747 ), .C(\U1/keyexpantion/SB0/n2746 ), .D(
        \U1/keyexpantion/SB0/n2745 ), .E(\U1/keyexpantion/SB0/n2744 ), .F(
        \U1/keyexpantion/SB0/n2743 ), .Y(\U1/keyexpantion/SB0/n2828 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U264  ( .A0(
        \U1/keyexpantion/SB0/n2940 ), .A1(\U1/keyexpantion/SB0/n2749 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .B1(\U1/keyexpantion/SB0/n2875 ), .Y(
        \U1/keyexpantion/SB0/n2750 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U263  ( .A0(
        \U1/keyexpantion/SB0/n2801 ), .A1(\U1/keyexpantion/SB0/n2967 ), .B0(
        \U1/keyexpantion/SB0/n2751 ), .B1(\U1/keyexpantion/SB0/n2957 ), .C0(
        \U1/keyexpantion/SB0/n2750 ), .Y(\U1/keyexpantion/SB0/n2763 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U262  ( .AN(
        \U1/keyexpantion/SB0/n2755 ), .B(\U1/keyexpantion/SB0/n2754 ), .C(
        \U1/keyexpantion/SB0/n2753 ), .D(\U1/keyexpantion/SB0/n2752 ), .Y(
        \U1/keyexpantion/SB0/n2762 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U261  ( .A0(
        \U1/keyexpantion/SB0/n2960 ), .A1(\U1/keyexpantion/SB0/n2756 ), .B0(
        \U1/keyexpantion/SB0/n2951 ), .Y(\U1/keyexpantion/SB0/n2760 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U260  ( .A(
        \U1/keyexpantion/SB0/n2927 ), .B(\U1/keyexpantion/SB0/n2932 ), .Y(
        \U1/keyexpantion/SB0/n2757 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U259  ( .A0(
        \U1/keyexpantion/SB0/n2882 ), .A1(\U1/keyexpantion/SB0/n2757 ), .B0(
        \U1/keyexpantion/SB0/n2883 ), .B1(\U1/keyexpantion/SB0/n2829 ), .Y(
        \U1/keyexpantion/SB0/n2758 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U258  ( .A(
        \U1/keyexpantion/SB0/n2760 ), .B(\U1/keyexpantion/SB0/n2759 ), .C(
        \U1/keyexpantion/SB0/n2758 ), .Y(\U1/keyexpantion/SB0/n2761 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U257  ( .A(\U1/keyexpantion/SB0/n2821 ), 
        .B(\U1/keyexpantion/SB0/n2869 ), .C(\U1/keyexpantion/SB0/n2828 ), .D(
        \U1/keyexpantion/SB0/n2763 ), .E(\U1/keyexpantion/SB0/n2762 ), .F(
        \U1/keyexpantion/SB0/n2761 ), .Y(\U1/keyexpantion/SB0/n2936 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U256  ( .A(\U1/keyexpantion/SB0/n2848 ), 
        .B(\U1/keyexpantion/SB0/n2893 ), .C(\U1/keyexpantion/SB0/n2797 ), .D(
        \U1/keyexpantion/SB0/n2936 ), .Y(\U1/keyexpantion/SB0/n2777 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U255  ( .A0(
        \U1/keyexpantion/SB0/n2916 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2764 ), .B1(\U1/keyexpantion/SB0/n2932 ), .Y(
        \U1/keyexpantion/SB0/n2765 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U254  ( .A0(
        \U1/keyexpantion/SB0/n2921 ), .A1(\U1/keyexpantion/SB0/n2939 ), .B0(
        \U1/keyexpantion/SB0/n2952 ), .B1(\U1/keyexpantion/SB0/n2960 ), .C0(
        \U1/keyexpantion/SB0/n2765 ), .Y(\U1/keyexpantion/SB0/n2776 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U253  ( .A(\U1/keyexpantion/SB0/n2766 ), 
        .Y(\U1/keyexpantion/SB0/n2769 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U252  ( .A0(
        \U1/keyexpantion/SB0/n2767 ), .A1(\U1/keyexpantion/SB0/n2872 ), .B0(
        \U1/keyexpantion/SB0/n2800 ), .B1(\U1/keyexpantion/SB0/n2852 ), .Y(
        \U1/keyexpantion/SB0/n2768 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U251  ( .A0(
        \U1/keyexpantion/SB0/n2940 ), .A1(\U1/keyexpantion/SB0/n2769 ), .B0(
        \U1/keyexpantion/SB0/n2922 ), .B1(\U1/keyexpantion/SB0/n2850 ), .C0(
        \U1/keyexpantion/SB0/n2768 ), .Y(\U1/keyexpantion/SB0/n2775 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U250  ( .A0(
        \U1/keyexpantion/SB0/n2962 ), .A1(\U1/keyexpantion/SB0/n2818 ), .B0(
        \U1/keyexpantion/SB0/n2942 ), .Y(\U1/keyexpantion/SB0/n2773 ) );
  AND4_X0P5M_A12TL \U1/keyexpantion/SB0/U249  ( .A(\U1/keyexpantion/SB0/n2773 ), .B(\U1/keyexpantion/SB0/n2772 ), .C(\U1/keyexpantion/SB0/n2771 ), .D(
        \U1/keyexpantion/SB0/n2770 ), .Y(\U1/keyexpantion/SB0/n2774 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U248  ( .AN(
        \U1/keyexpantion/SB0/n2777 ), .B(\U1/keyexpantion/SB0/n2776 ), .C(
        \U1/keyexpantion/SB0/n2775 ), .D(\U1/keyexpantion/SB0/n2774 ), .Y(
        \U1/keyexpantion/ws [27]) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U247  ( .A0(
        \U1/keyexpantion/SB0/n2792 ), .A1(\U1/keyexpantion/SB0/n2928 ), .B0(
        \U1/keyexpantion/SB0/n2851 ), .Y(\U1/keyexpantion/SB0/n2789 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U246  ( .A(
        \U1/keyexpantion/SB0/n2780 ), .B(\U1/keyexpantion/SB0/n2779 ), .C(
        \U1/keyexpantion/SB0/n2778 ), .Y(\U1/keyexpantion/SB0/n2788 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U245  ( .A(\U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2951 ), .Y(\U1/keyexpantion/SB0/n2783 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U244  ( .A(\U1/keyexpantion/SB0/n2922 ), .B(\U1/keyexpantion/SB0/n2835 ), .Y(\U1/keyexpantion/SB0/n2781 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U243  ( .A0(
        \U1/keyexpantion/SB0/n2783 ), .A1(\U1/keyexpantion/SB0/n2782 ), .B0(
        \U1/keyexpantion/SB0/n2781 ), .B1(\U1/keyexpantion/SB0/n2945 ), .C0(
        \U1/keyexpantion/SB0/n2928 ), .C1(\U1/keyexpantion/SB0/n2833 ), .Y(
        \U1/keyexpantion/SB0/n2787 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U242  ( .A0(
        \U1/keyexpantion/SB0/n2884 ), .A1(\U1/keyexpantion/SB0/n2785 ), .B0(
        \U1/keyexpantion/SB0/n2967 ), .B1(\U1/keyexpantion/SB0/n2957 ), .C0(
        \U1/keyexpantion/SB0/n2930 ), .C1(\U1/keyexpantion/SB0/n2784 ), .Y(
        \U1/keyexpantion/SB0/n2786 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U241  ( .A(\U1/keyexpantion/SB0/n2791 ), 
        .B(\U1/keyexpantion/SB0/n2790 ), .C(\U1/keyexpantion/SB0/n2789 ), .D(
        \U1/keyexpantion/SB0/n2788 ), .E(\U1/keyexpantion/SB0/n2787 ), .F(
        \U1/keyexpantion/SB0/n2786 ), .Y(\U1/keyexpantion/SB0/n2937 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U240  ( .A0(
        \U1/keyexpantion/SB0/n2792 ), .A1(\U1/keyexpantion/SB0/n2801 ), .B0(
        \U1/keyexpantion/SB0/n2872 ), .Y(\U1/keyexpantion/SB0/n2827 ) );
  AOI31_X0P5M_A12TL \U1/keyexpantion/SB0/U239  ( .A0(
        \U1/keyexpantion/SB0/n2917 ), .A1(\U1/keyexpantion/SB0/n2930 ), .A2(
        \U1/keyexpantion/SB0/n2849 ), .B0(\U1/keyexpantion/SB0/n2946 ), .Y(
        \U1/keyexpantion/SB0/n2826 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U238  ( .A(
        \U1/keyexpantion/SB0/n2796 ), .B(\U1/keyexpantion/SB0/n2795 ), .C(
        \U1/keyexpantion/SB0/n2794 ), .D(\U1/keyexpantion/SB0/n2793 ), .Y(
        \U1/keyexpantion/SB0/n2823 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U237  ( .A(\U1/keyexpantion/SB0/n2797 ), 
        .Y(\U1/keyexpantion/SB0/n2820 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U236  ( .A(\U1/keyexpantion/SB0/n2798 ), 
        .Y(\U1/keyexpantion/SB0/n2814 ) );
  OAI21B_X0P5M_A12TL \U1/keyexpantion/SB0/U235  ( .A0(
        \U1/keyexpantion/SB0/n2800 ), .A1(\U1/keyexpantion/SB0/n2958 ), .B0N(
        \U1/keyexpantion/SB0/n2799 ), .Y(\U1/keyexpantion/SB0/n2813 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U234  ( .A0(
        \U1/keyexpantion/SB0/n2965 ), .A1(\U1/keyexpantion/SB0/n2801 ), .B0(
        \U1/keyexpantion/SB0/n2851 ), .B1(\U1/keyexpantion/SB0/n2932 ), .C0(
        \U1/keyexpantion/SB0/n2946 ), .C1(\U1/keyexpantion/SB0/n2967 ), .Y(
        \U1/keyexpantion/SB0/n2812 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U233  ( .AN(
        \U1/keyexpantion/SB0/n2805 ), .B(\U1/keyexpantion/SB0/n2804 ), .C(
        \U1/keyexpantion/SB0/n2803 ), .D(\U1/keyexpantion/SB0/n2802 ), .Y(
        \U1/keyexpantion/SB0/n2811 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U232  ( .A(
        \U1/keyexpantion/SB0/n2809 ), .B(\U1/keyexpantion/SB0/n2808 ), .C(
        \U1/keyexpantion/SB0/n2807 ), .D(\U1/keyexpantion/SB0/n2806 ), .Y(
        \U1/keyexpantion/SB0/n2810 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U231  ( .A(\U1/keyexpantion/SB0/n2815 ), 
        .B(\U1/keyexpantion/SB0/n2814 ), .C(\U1/keyexpantion/SB0/n2813 ), .D(
        \U1/keyexpantion/SB0/n2812 ), .E(\U1/keyexpantion/SB0/n2811 ), .F(
        \U1/keyexpantion/SB0/n2810 ), .Y(\U1/keyexpantion/SB0/n2816 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U230  ( .A(\U1/keyexpantion/SB0/n2816 ), 
        .Y(\U1/keyexpantion/SB0/n2915 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U229  ( .A0(
        \U1/keyexpantion/SB0/n2884 ), .A1(\U1/keyexpantion/SB0/n2927 ), .B0(
        \U1/keyexpantion/SB0/n2967 ), .B1(\U1/keyexpantion/SB0/n2966 ), .Y(
        \U1/keyexpantion/SB0/n2817 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U228  ( .A0(
        \U1/keyexpantion/SB0/n2874 ), .A1(\U1/keyexpantion/SB0/n2818 ), .B0(
        \U1/keyexpantion/SB0/n2919 ), .B1(\U1/keyexpantion/SB0/n2941 ), .C0(
        \U1/keyexpantion/SB0/n2817 ), .Y(\U1/keyexpantion/SB0/n2819 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U227  ( .AN(
        \U1/keyexpantion/SB0/n2821 ), .B(\U1/keyexpantion/SB0/n2820 ), .C(
        \U1/keyexpantion/SB0/n2915 ), .D(\U1/keyexpantion/SB0/n2819 ), .Y(
        \U1/keyexpantion/SB0/n2822 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U226  ( .A(\U1/keyexpantion/SB0/n2827 ), 
        .B(\U1/keyexpantion/SB0/n2826 ), .C(\U1/keyexpantion/SB0/n2825 ), .D(
        \U1/keyexpantion/SB0/n2824 ), .E(\U1/keyexpantion/SB0/n2823 ), .F(
        \U1/keyexpantion/SB0/n2822 ), .Y(\U1/keyexpantion/SB0/n2892 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U225  ( .A(\U1/keyexpantion/SB0/n2828 ), 
        .Y(\U1/keyexpantion/SB0/n2832 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U224  ( .A0(
        \U1/keyexpantion/SB0/n2830 ), .A1(\U1/keyexpantion/SB0/n2829 ), .B0(
        \U1/keyexpantion/SB0/n2876 ), .B1(\U1/keyexpantion/SB0/n2835 ), .Y(
        \U1/keyexpantion/SB0/n2831 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U223  ( .A0(
        \U1/keyexpantion/SB0/n2946 ), .A1(\U1/keyexpantion/SB0/n2833 ), .B0(
        \U1/keyexpantion/SB0/n2832 ), .C0(\U1/keyexpantion/SB0/n2831 ), .Y(
        \U1/keyexpantion/SB0/n2847 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U222  ( .A0(
        \U1/keyexpantion/SB0/n2834 ), .A1(\U1/keyexpantion/SB0/n2918 ), .B0(
        \U1/keyexpantion/SB0/n2947 ), .Y(\U1/keyexpantion/SB0/n2839 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U221  ( .A0(
        \U1/keyexpantion/SB0/n2835 ), .A1(\U1/keyexpantion/SB0/n2921 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2838 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U220  ( .A(
        \U1/keyexpantion/SB0/n2839 ), .B(\U1/keyexpantion/SB0/n2838 ), .C(
        \U1/keyexpantion/SB0/n2837 ), .D(\U1/keyexpantion/SB0/n2836 ), .Y(
        \U1/keyexpantion/SB0/n2846 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U219  ( .A(\U1/keyexpantion/SB0/n2877 ), .B(\U1/keyexpantion/SB0/n2840 ), .Y(\U1/keyexpantion/SB0/n2844 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U218  ( .A(\U1/keyexpantion/SB0/n2841 ), .B(\U1/keyexpantion/SB0/n2882 ), .Y(\U1/keyexpantion/SB0/n2843 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U217  ( .A0(
        \U1/keyexpantion/SB0/n2844 ), .A1(\U1/keyexpantion/SB0/n2964 ), .B0(
        \U1/keyexpantion/SB0/n2843 ), .B1(\U1/keyexpantion/SB0/n2928 ), .C0(
        \U1/keyexpantion/SB0/n2842 ), .C1(\U1/keyexpantion/SB0/n2929 ), .Y(
        \U1/keyexpantion/SB0/n2845 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U216  ( .A(\U1/keyexpantion/SB0/n2937 ), 
        .B(\U1/keyexpantion/SB0/n2892 ), .C(\U1/keyexpantion/SB0/n2848 ), .D(
        \U1/keyexpantion/SB0/n2847 ), .E(\U1/keyexpantion/SB0/n2846 ), .F(
        \U1/keyexpantion/SB0/n2845 ), .Y(\U1/keyexpantion/ws [28]) );
  AOI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U215  ( .A1N(
        \U1/keyexpantion/SB0/n2850 ), .A0(\U1/keyexpantion/SB0/n2849 ), .B0(
        \U1/keyexpantion/SB0/n2927 ), .Y(\U1/keyexpantion/SB0/n2866 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U214  ( .A(\U1/keyexpantion/SB0/n2940 ), .B(\U1/keyexpantion/SB0/n2921 ), .Y(\U1/keyexpantion/SB0/n2853 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U213  ( .A0(
        \U1/keyexpantion/SB0/n2964 ), .A1(\U1/keyexpantion/SB0/n2854 ), .B0(
        \U1/keyexpantion/SB0/n2853 ), .B1(\U1/keyexpantion/SB0/n2967 ), .C0(
        \U1/keyexpantion/SB0/n2852 ), .C1(\U1/keyexpantion/SB0/n2851 ), .Y(
        \U1/keyexpantion/SB0/n2865 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U212  ( .A(\U1/keyexpantion/SB0/n2855 ), 
        .Y(\U1/keyexpantion/SB0/n2858 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U211  ( .AN(
        \U1/keyexpantion/SB0/n2859 ), .B(\U1/keyexpantion/SB0/n2858 ), .C(
        \U1/keyexpantion/SB0/n2857 ), .D(\U1/keyexpantion/SB0/n2856 ), .Y(
        \U1/keyexpantion/SB0/n2864 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U210  ( .A(
        \U1/keyexpantion/SB0/n2862 ), .B(\U1/keyexpantion/SB0/n2861 ), .C(
        \U1/keyexpantion/SB0/n2860 ), .Y(\U1/keyexpantion/SB0/n2863 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U209  ( .A(\U1/keyexpantion/SB0/n2868 ), 
        .B(\U1/keyexpantion/SB0/n2867 ), .C(\U1/keyexpantion/SB0/n2866 ), .D(
        \U1/keyexpantion/SB0/n2865 ), .E(\U1/keyexpantion/SB0/n2864 ), .F(
        \U1/keyexpantion/SB0/n2863 ), .Y(\U1/keyexpantion/SB0/n2938 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U208  ( .A(\U1/keyexpantion/SB0/n2869 ), 
        .Y(\U1/keyexpantion/SB0/n2871 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U207  ( .A0(
        \U1/keyexpantion/SB0/n2951 ), .A1(\U1/keyexpantion/SB0/n2948 ), .B0(
        \U1/keyexpantion/SB0/n2952 ), .B1(\U1/keyexpantion/SB0/n2950 ), .Y(
        \U1/keyexpantion/SB0/n2870 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U206  ( .A0(
        \U1/keyexpantion/SB0/n2927 ), .A1(\U1/keyexpantion/SB0/n2872 ), .B0(
        \U1/keyexpantion/SB0/n2871 ), .C0(\U1/keyexpantion/SB0/n2870 ), .Y(
        \U1/keyexpantion/SB0/n2891 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U205  ( .A0(
        \U1/keyexpantion/SB0/n2874 ), .A1(\U1/keyexpantion/SB0/n2951 ), .B0(
        \U1/keyexpantion/SB0/n2873 ), .Y(\U1/keyexpantion/SB0/n2880 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U204  ( .A0(
        \U1/keyexpantion/SB0/n2877 ), .A1(\U1/keyexpantion/SB0/n2876 ), .B0(
        \U1/keyexpantion/SB0/n2875 ), .Y(\U1/keyexpantion/SB0/n2879 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U203  ( .AN(
        \U1/keyexpantion/SB0/n2881 ), .B(\U1/keyexpantion/SB0/n2880 ), .C(
        \U1/keyexpantion/SB0/n2879 ), .D(\U1/keyexpantion/SB0/n2878 ), .Y(
        \U1/keyexpantion/SB0/n2890 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U202  ( .A0(
        \U1/keyexpantion/SB0/n2947 ), .A1(\U1/keyexpantion/SB0/n2883 ), .B0(
        \U1/keyexpantion/SB0/n2882 ), .Y(\U1/keyexpantion/SB0/n2887 ) );
  OA22_X0P5M_A12TL \U1/keyexpantion/SB0/U201  ( .A0(
        \U1/keyexpantion/SB0/n2929 ), .A1(\U1/keyexpantion/SB0/n2885 ), .B0(
        \U1/keyexpantion/SB0/n2966 ), .B1(\U1/keyexpantion/SB0/n2884 ), .Y(
        \U1/keyexpantion/SB0/n2886 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U200  ( .A0(
        \U1/keyexpantion/SB0/n2888 ), .A1(\U1/keyexpantion/SB0/n2928 ), .B0(
        \U1/keyexpantion/SB0/n2887 ), .C0(\U1/keyexpantion/SB0/n2886 ), .Y(
        \U1/keyexpantion/SB0/n2889 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U199  ( .A(\U1/keyexpantion/SB0/n2938 ), 
        .B(\U1/keyexpantion/SB0/n2893 ), .C(\U1/keyexpantion/SB0/n2892 ), .D(
        \U1/keyexpantion/SB0/n2891 ), .E(\U1/keyexpantion/SB0/n2890 ), .F(
        \U1/keyexpantion/SB0/n2889 ), .Y(\U1/keyexpantion/ws [29]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U198  ( .A0(
        \U1/keyexpantion/SB0/n3221 ), .A1(\U1/keyexpantion/SB0/n3241 ), .B0(
        \U1/keyexpantion/SB0/n3262 ), .B1(\U1/keyexpantion/SB0/n3252 ), .Y(
        \U1/keyexpantion/SB0/n2894 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U197  ( .A0(
        \U1/keyexpantion/SB0/n3172 ), .A1(\U1/keyexpantion/SB0/n3266 ), .B0(
        \U1/keyexpantion/SB0/n3122 ), .B1(\U1/keyexpantion/SB0/n3193 ), .C0(
        \U1/keyexpantion/SB0/n2894 ), .Y(\U1/keyexpantion/SB0/n2900 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U196  ( .A(
        \U1/keyexpantion/SB0/n3247 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3056 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U195  ( .A(
        \U1/keyexpantion/SB0/n3221 ), .B(\U1/keyexpantion/SB0/n3197 ), .Y(
        \U1/keyexpantion/SB0/n3037 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U194  ( .A(
        \U1/keyexpantion/SB0/n3241 ), .B(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3005 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U193  ( .A(
        \U1/keyexpantion/SB0/n3161 ), .B(\U1/keyexpantion/SB0/n3204 ), .Y(
        \U1/keyexpantion/SB0/n3024 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U192  ( .A(
        \U1/keyexpantion/SB0/n3056 ), .B(\U1/keyexpantion/SB0/n3037 ), .C(
        \U1/keyexpantion/SB0/n3005 ), .D(\U1/keyexpantion/SB0/n3024 ), .Y(
        \U1/keyexpantion/SB0/n2899 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U191  ( .A(
        \U1/keyexpantion/SB0/n3267 ), .B(\U1/keyexpantion/SB0/n3245 ), .Y(
        \U1/keyexpantion/SB0/n3150 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U190  ( .A0(
        \U1/keyexpantion/SB0/n3198 ), .A1(\U1/keyexpantion/SB0/n3150 ), .B0(
        \U1/keyexpantion/SB0/n3251 ), .Y(\U1/keyexpantion/SB0/n2897 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U189  ( .A0(
        \U1/keyexpantion/SB0/n3248 ), .A1(\U1/keyexpantion/SB0/n3139 ), .B0(
        \U1/keyexpantion/SB0/n3151 ), .Y(\U1/keyexpantion/SB0/n2896 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U188  ( .A0(
        \U1/keyexpantion/SB0/n3156 ), .A1(\U1/keyexpantion/SB0/n3196 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n2895 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U187  ( .A(
        \U1/keyexpantion/SB0/n3240 ), .B(\U1/keyexpantion/SB0/n3248 ), .Y(
        \U1/keyexpantion/SB0/n3123 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U186  ( .A(
        \U1/keyexpantion/SB0/n2897 ), .B(\U1/keyexpantion/SB0/n2896 ), .C(
        \U1/keyexpantion/SB0/n2895 ), .D(\U1/keyexpantion/SB0/n3123 ), .Y(
        \U1/keyexpantion/SB0/n2898 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U185  ( .A(\U1/keyexpantion/SB0/n2903 ), 
        .B(\U1/keyexpantion/SB0/n2902 ), .C(\U1/keyexpantion/SB0/n2901 ), .D(
        \U1/keyexpantion/SB0/n2900 ), .E(\U1/keyexpantion/SB0/n2899 ), .F(
        \U1/keyexpantion/SB0/n2898 ), .Y(\U1/keyexpantion/SB0/n3271 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U184  ( .A0(
        \U1/keyexpantion/SB0/n3077 ), .A1(\U1/keyexpantion/SB0/n3252 ), .B0(
        \U1/keyexpantion/SB0/n3260 ), .B1(\U1/keyexpantion/SB0/n3195 ), .C0(
        \U1/keyexpantion/SB0/n3271 ), .Y(\U1/keyexpantion/SB0/n2904 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U183  ( .A(\U1/keyexpantion/SB0/n2904 ), 
        .Y(\U1/keyexpantion/SB0/n2911 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U182  ( .A(\U1/keyexpantion/SB0/n3204 ), .B(\U1/keyexpantion/SB0/n2991 ), .Y(\U1/keyexpantion/SB0/n3113 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U181  ( .A1N(
        \U1/keyexpantion/SB0/n3113 ), .A0(\U1/keyexpantion/SB0/n3222 ), .B0(
        \U1/keyexpantion/SB0/n3194 ), .Y(\U1/keyexpantion/SB0/n2907 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U180  ( .A0(
        \U1/keyexpantion/SB0/n3162 ), .A1(\U1/keyexpantion/SB0/n3070 ), .B0(
        \U1/keyexpantion/SB0/n3221 ), .Y(\U1/keyexpantion/SB0/n2906 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U179  ( .A0(
        \U1/keyexpantion/SB0/n3248 ), .A1(\U1/keyexpantion/SB0/n3203 ), .B0(
        \U1/keyexpantion/SB0/n3242 ), .Y(\U1/keyexpantion/SB0/n2905 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U178  ( .A(
        \U1/keyexpantion/SB0/n3219 ), .B(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3020 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U177  ( .A(
        \U1/keyexpantion/SB0/n2907 ), .B(\U1/keyexpantion/SB0/n2906 ), .C(
        \U1/keyexpantion/SB0/n2905 ), .D(\U1/keyexpantion/SB0/n3020 ), .Y(
        \U1/keyexpantion/SB0/n2910 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U176  ( .A(\U1/keyexpantion/SB0/n3218 ), .B(\U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n3249 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U175  ( .A(\U1/keyexpantion/SB0/n3240 ), .B(\U1/keyexpantion/SB0/n3196 ), .Y(\U1/keyexpantion/SB0/n2908 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U174  ( .A0(
        \U1/keyexpantion/SB0/n3249 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n2908 ), .B1(\U1/keyexpantion/SB0/n3230 ), .C0(
        \U1/keyexpantion/SB0/n3173 ), .C1(\U1/keyexpantion/SB0/n3175 ), .Y(
        \U1/keyexpantion/SB0/n2909 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U173  ( .A(\U1/keyexpantion/SB0/n2914 ), 
        .B(\U1/keyexpantion/SB0/n2913 ), .C(\U1/keyexpantion/SB0/n2912 ), .D(
        \U1/keyexpantion/SB0/n2911 ), .E(\U1/keyexpantion/SB0/n2910 ), .F(
        \U1/keyexpantion/SB0/n2909 ), .Y(\U1/keyexpantion/ws [2]) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U172  ( .A0(
        \U1/keyexpantion/SB0/n2917 ), .A1(\U1/keyexpantion/SB0/n2957 ), .B0(
        \U1/keyexpantion/SB0/n2916 ), .B1(\U1/keyexpantion/SB0/n2964 ), .C0(
        \U1/keyexpantion/SB0/n2915 ), .Y(\U1/keyexpantion/SB0/n2935 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U171  ( .A0(
        \U1/keyexpantion/SB0/n2918 ), .A1(\U1/keyexpantion/SB0/n2962 ), .B0(
        \U1/keyexpantion/SB0/n2951 ), .Y(\U1/keyexpantion/SB0/n2926 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U170  ( .A0(
        \U1/keyexpantion/SB0/n2942 ), .A1(\U1/keyexpantion/SB0/n2919 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2925 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U169  ( .A0(
        \U1/keyexpantion/SB0/n2922 ), .A1(\U1/keyexpantion/SB0/n2921 ), .B0(
        \U1/keyexpantion/SB0/n2920 ), .Y(\U1/keyexpantion/SB0/n2924 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U168  ( .A(
        \U1/keyexpantion/SB0/n2926 ), .B(\U1/keyexpantion/SB0/n2925 ), .C(
        \U1/keyexpantion/SB0/n2924 ), .D(\U1/keyexpantion/SB0/n2923 ), .Y(
        \U1/keyexpantion/SB0/n2934 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U167  ( .A(
        \U1/keyexpantion/SB0/n2957 ), .B(\U1/keyexpantion/SB0/n2927 ), .Y(
        \U1/keyexpantion/SB0/n2959 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U166  ( .A(\U1/keyexpantion/SB0/n2947 ), .B(\U1/keyexpantion/SB0/n2959 ), .Y(\U1/keyexpantion/SB0/n2931 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U165  ( .A0(
        \U1/keyexpantion/SB0/n2945 ), .A1(\U1/keyexpantion/SB0/n2932 ), .B0(
        \U1/keyexpantion/SB0/n2931 ), .B1(\U1/keyexpantion/SB0/n2930 ), .C0(
        \U1/keyexpantion/SB0/n2929 ), .C1(\U1/keyexpantion/SB0/n2928 ), .Y(
        \U1/keyexpantion/SB0/n2933 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U164  ( .A(\U1/keyexpantion/SB0/n2938 ), 
        .B(\U1/keyexpantion/SB0/n2937 ), .C(\U1/keyexpantion/SB0/n2936 ), .D(
        \U1/keyexpantion/SB0/n2935 ), .E(\U1/keyexpantion/SB0/n2934 ), .F(
        \U1/keyexpantion/SB0/n2933 ), .Y(\U1/keyexpantion/ws [30]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U163  ( .A0(
        \U1/keyexpantion/SB0/n2942 ), .A1(\U1/keyexpantion/SB0/n2941 ), .B0(
        \U1/keyexpantion/SB0/n2940 ), .B1(\U1/keyexpantion/SB0/n2939 ), .Y(
        \U1/keyexpantion/SB0/n2943 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U162  ( .A0(
        \U1/keyexpantion/SB0/n2946 ), .A1(\U1/keyexpantion/SB0/n2945 ), .B0(
        \U1/keyexpantion/SB0/n2944 ), .C0(\U1/keyexpantion/SB0/n2943 ), .Y(
        \U1/keyexpantion/SB0/n2970 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U161  ( .A1N(
        \U1/keyexpantion/SB0/n2949 ), .A0(\U1/keyexpantion/SB0/n2948 ), .B0(
        \U1/keyexpantion/SB0/n2947 ), .Y(\U1/keyexpantion/SB0/n2956 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U160  ( .A0(
        \U1/keyexpantion/SB0/n2952 ), .A1(\U1/keyexpantion/SB0/n2951 ), .B0(
        \U1/keyexpantion/SB0/n2950 ), .Y(\U1/keyexpantion/SB0/n2955 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U159  ( .A(
        \U1/keyexpantion/SB0/n2956 ), .B(\U1/keyexpantion/SB0/n2955 ), .C(
        \U1/keyexpantion/SB0/n2954 ), .D(\U1/keyexpantion/SB0/n2953 ), .Y(
        \U1/keyexpantion/SB0/n2969 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U158  ( .A(
        \U1/keyexpantion/SB0/n2958 ), .B(\U1/keyexpantion/SB0/n2957 ), .Y(
        \U1/keyexpantion/SB0/n2961 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U157  ( .A0(
        \U1/keyexpantion/SB0/n2962 ), .A1(\U1/keyexpantion/SB0/n2961 ), .B0(
        \U1/keyexpantion/SB0/n2960 ), .B1(\U1/keyexpantion/SB0/n2959 ), .Y(
        \U1/keyexpantion/SB0/n2963 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U156  ( .A0(
        \U1/keyexpantion/SB0/n2967 ), .A1(\U1/keyexpantion/SB0/n2966 ), .B0(
        \U1/keyexpantion/SB0/n2965 ), .B1(\U1/keyexpantion/SB0/n2964 ), .C0(
        \U1/keyexpantion/SB0/n2963 ), .Y(\U1/keyexpantion/SB0/n2968 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U155  ( .A(\U1/keyexpantion/SB0/n2973 ), 
        .B(\U1/keyexpantion/SB0/n2972 ), .C(\U1/keyexpantion/SB0/n2971 ), .D(
        \U1/keyexpantion/SB0/n2970 ), .E(\U1/keyexpantion/SB0/n2969 ), .F(
        \U1/keyexpantion/SB0/n2968 ), .Y(\U1/keyexpantion/ws [31]) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U154  ( .A(
        \U1/keyexpantion/SB0/n3077 ), .B(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3254 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U153  ( .AN(
        \U1/keyexpantion/SB0/n2976 ), .B(\U1/keyexpantion/SB0/n2975 ), .C(
        \U1/keyexpantion/SB0/n2974 ), .D(\U1/keyexpantion/SB0/n3254 ), .Y(
        \U1/keyexpantion/SB0/n2983 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U152  ( .A0(
        \U1/keyexpantion/SB0/n2977 ), .A1(\U1/keyexpantion/SB0/n3221 ), .B0(
        \U1/keyexpantion/SB0/n3139 ), .Y(\U1/keyexpantion/SB0/n2979 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U149  ( .A(\U1/keyexpantion/SB0/n3195 ), .B(\U1/keyexpantion/SB0/n3242 ), .Y(\U1/keyexpantion/SB0/n3206 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U148  ( .A0(
        \U1/keyexpantion/SB0/n3085 ), .A1(\U1/keyexpantion/SB0/n3264 ), .B0(
        \U1/keyexpantion/SB0/n3206 ), .B1(\U1/keyexpantion/SB0/n3217 ), .C0(
        \U1/keyexpantion/SB0/n3258 ), .C1(\U1/keyexpantion/SB0/n3267 ), .Y(
        \U1/keyexpantion/SB0/n2981 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U147  ( .A(\U1/keyexpantion/SB0/n2986 ), 
        .B(\U1/keyexpantion/SB0/n2985 ), .C(\U1/keyexpantion/SB0/n2984 ), .D(
        \U1/keyexpantion/SB0/n2983 ), .E(\U1/keyexpantion/SB0/n2982 ), .F(
        \U1/keyexpantion/SB0/n2981 ), .Y(\U1/keyexpantion/SB0/n3169 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U146  ( .AN(
        \U1/keyexpantion/SB0/n2990 ), .B(\U1/keyexpantion/SB0/n2989 ), .C(
        \U1/keyexpantion/SB0/n2988 ), .D(\U1/keyexpantion/SB0/n2987 ), .Y(
        \U1/keyexpantion/SB0/n3000 ) );
  AOI222_X0P5M_A12TL \U1/keyexpantion/SB0/U145  ( .A0(
        \U1/keyexpantion/SB0/n3252 ), .A1(\U1/keyexpantion/SB0/n3162 ), .B0(
        \U1/keyexpantion/SB0/n3247 ), .B1(\U1/keyexpantion/SB0/n3161 ), .C0(
        \U1/keyexpantion/SB0/n2991 ), .C1(\U1/keyexpantion/SB0/n3262 ), .Y(
        \U1/keyexpantion/SB0/n2999 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U144  ( .A0(
        \U1/keyexpantion/SB0/n3216 ), .A1(\U1/keyexpantion/SB0/n3122 ), .B0(
        \U1/keyexpantion/SB0/n2992 ), .B1(\U1/keyexpantion/SB0/n3085 ), .Y(
        \U1/keyexpantion/SB0/n2993 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U143  ( .A0(
        \U1/keyexpantion/SB0/n3139 ), .A1(\U1/keyexpantion/SB0/n3156 ), .B0(
        \U1/keyexpantion/SB0/n3155 ), .B1(\U1/keyexpantion/SB0/n3219 ), .C0(
        \U1/keyexpantion/SB0/n2993 ), .Y(\U1/keyexpantion/SB0/n2998 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U142  ( .A(
        \U1/keyexpantion/SB0/n3227 ), .B(\U1/keyexpantion/SB0/n3266 ), .Y(
        \U1/keyexpantion/SB0/n2995 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U141  ( .A0(
        \U1/keyexpantion/SB0/n3077 ), .A1(\U1/keyexpantion/SB0/n2996 ), .B0(
        \U1/keyexpantion/SB0/n3248 ), .B1(\U1/keyexpantion/SB0/n2995 ), .C0(
        \U1/keyexpantion/SB0/n2994 ), .Y(\U1/keyexpantion/SB0/n2997 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U140  ( .AN(
        \U1/keyexpantion/SB0/n3000 ), .B(\U1/keyexpantion/SB0/n2999 ), .C(
        \U1/keyexpantion/SB0/n2998 ), .D(\U1/keyexpantion/SB0/n2997 ), .Y(
        \U1/keyexpantion/SB0/n3214 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U139  ( .A(\U1/keyexpantion/SB0/n3001 ), 
        .Y(\U1/keyexpantion/SB0/n3017 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U138  ( .A0(
        \U1/keyexpantion/SB0/n3106 ), .A1(\U1/keyexpantion/SB0/n3175 ), .B0(
        \U1/keyexpantion/SB0/n3002 ), .Y(\U1/keyexpantion/SB0/n3016 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U137  ( .A0(
        \U1/keyexpantion/SB0/n3248 ), .A1(\U1/keyexpantion/SB0/n3247 ), .B0(
        \U1/keyexpantion/SB0/n3218 ), .B1(\U1/keyexpantion/SB0/n3003 ), .Y(
        \U1/keyexpantion/SB0/n3004 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U136  ( .A0(
        \U1/keyexpantion/SB0/n3229 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n3245 ), .B1(\U1/keyexpantion/SB0/n3257 ), .C0(
        \U1/keyexpantion/SB0/n3004 ), .Y(\U1/keyexpantion/SB0/n3015 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U135  ( .A(
        \U1/keyexpantion/SB0/n3008 ), .B(\U1/keyexpantion/SB0/n3007 ), .C(
        \U1/keyexpantion/SB0/n3006 ), .D(\U1/keyexpantion/SB0/n3005 ), .Y(
        \U1/keyexpantion/SB0/n3014 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U134  ( .AN(
        \U1/keyexpantion/SB0/n3012 ), .B(\U1/keyexpantion/SB0/n3011 ), .C(
        \U1/keyexpantion/SB0/n3010 ), .D(\U1/keyexpantion/SB0/n3009 ), .Y(
        \U1/keyexpantion/SB0/n3013 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U133  ( .A(\U1/keyexpantion/SB0/n3018 ), 
        .B(\U1/keyexpantion/SB0/n3017 ), .C(\U1/keyexpantion/SB0/n3016 ), .D(
        \U1/keyexpantion/SB0/n3015 ), .E(\U1/keyexpantion/SB0/n3014 ), .F(
        \U1/keyexpantion/SB0/n3013 ), .Y(\U1/keyexpantion/SB0/n3118 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U132  ( .A0(
        \U1/keyexpantion/SB0/n3205 ), .A1(\U1/keyexpantion/SB0/n3122 ), .B0(
        \U1/keyexpantion/SB0/n3019 ), .Y(\U1/keyexpantion/SB0/n3034 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U131  ( .AN(
        \U1/keyexpantion/SB0/n3023 ), .B(\U1/keyexpantion/SB0/n3022 ), .C(
        \U1/keyexpantion/SB0/n3021 ), .D(\U1/keyexpantion/SB0/n3020 ), .Y(
        \U1/keyexpantion/SB0/n3033 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U130  ( .A(
        \U1/keyexpantion/SB0/n3239 ), .B(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3253 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U129  ( .A(
        \U1/keyexpantion/SB0/n3026 ), .B(\U1/keyexpantion/SB0/n3025 ), .C(
        \U1/keyexpantion/SB0/n3024 ), .D(\U1/keyexpantion/SB0/n3253 ), .Y(
        \U1/keyexpantion/SB0/n3032 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U128  ( .A(
        \U1/keyexpantion/SB0/n3030 ), .B(\U1/keyexpantion/SB0/n3029 ), .C(
        \U1/keyexpantion/SB0/n3028 ), .D(\U1/keyexpantion/SB0/n3027 ), .Y(
        \U1/keyexpantion/SB0/n3031 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U127  ( .A(\U1/keyexpantion/SB0/n3036 ), 
        .B(\U1/keyexpantion/SB0/n3035 ), .C(\U1/keyexpantion/SB0/n3034 ), .D(
        \U1/keyexpantion/SB0/n3033 ), .E(\U1/keyexpantion/SB0/n3032 ), .F(
        \U1/keyexpantion/SB0/n3031 ), .Y(\U1/keyexpantion/SB0/n3142 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U126  ( .AN(
        \U1/keyexpantion/SB0/n3040 ), .B(\U1/keyexpantion/SB0/n3039 ), .C(
        \U1/keyexpantion/SB0/n3038 ), .D(\U1/keyexpantion/SB0/n3037 ), .Y(
        \U1/keyexpantion/SB0/n3049 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U125  ( .A(
        \U1/keyexpantion/SB0/n3044 ), .B(\U1/keyexpantion/SB0/n3043 ), .C(
        \U1/keyexpantion/SB0/n3042 ), .D(\U1/keyexpantion/SB0/n3041 ), .Y(
        \U1/keyexpantion/SB0/n3048 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U124  ( .A(\U1/keyexpantion/SB0/n3204 ), .B(\U1/keyexpantion/SB0/n3240 ), .C(\U1/keyexpantion/SB0/n3242 ), .Y(
        \U1/keyexpantion/SB0/n3046 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U123  ( .A0(
        \U1/keyexpantion/SB0/n3046 ), .A1(\U1/keyexpantion/SB0/n3230 ), .B0(
        \U1/keyexpantion/SB0/n3085 ), .B1(\U1/keyexpantion/SB0/n3266 ), .C0(
        \U1/keyexpantion/SB0/n3045 ), .Y(\U1/keyexpantion/SB0/n3047 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U122  ( .A(\U1/keyexpantion/SB0/n3052 ), 
        .B(\U1/keyexpantion/SB0/n3051 ), .C(\U1/keyexpantion/SB0/n3050 ), .D(
        \U1/keyexpantion/SB0/n3049 ), .E(\U1/keyexpantion/SB0/n3048 ), .F(
        \U1/keyexpantion/SB0/n3047 ), .Y(\U1/keyexpantion/SB0/n3190 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U121  ( .A0(
        \U1/keyexpantion/SB0/n3085 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n3053 ), .Y(\U1/keyexpantion/SB0/n3067 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U120  ( .A0(
        \U1/keyexpantion/SB0/n3194 ), .A1(\U1/keyexpantion/SB0/n3196 ), .B0(
        \U1/keyexpantion/SB0/n3251 ), .B1(\U1/keyexpantion/SB0/n3161 ), .Y(
        \U1/keyexpantion/SB0/n3054 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U119  ( .A0(
        \U1/keyexpantion/SB0/n3105 ), .A1(\U1/keyexpantion/SB0/n3193 ), .B0(
        \U1/keyexpantion/SB0/n3106 ), .B1(\U1/keyexpantion/SB0/n3170 ), .C0(
        \U1/keyexpantion/SB0/n3054 ), .Y(\U1/keyexpantion/SB0/n3066 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U118  ( .A(\U1/keyexpantion/SB0/n3055 ), 
        .Y(\U1/keyexpantion/SB0/n3058 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U117  ( .AN(
        \U1/keyexpantion/SB0/n3059 ), .B(\U1/keyexpantion/SB0/n3058 ), .C(
        \U1/keyexpantion/SB0/n3057 ), .D(\U1/keyexpantion/SB0/n3056 ), .Y(
        \U1/keyexpantion/SB0/n3065 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U116  ( .A(
        \U1/keyexpantion/SB0/n3063 ), .B(\U1/keyexpantion/SB0/n3062 ), .C(
        \U1/keyexpantion/SB0/n3061 ), .D(\U1/keyexpantion/SB0/n3060 ), .Y(
        \U1/keyexpantion/SB0/n3064 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U115  ( .A(\U1/keyexpantion/SB0/n3069 ), 
        .B(\U1/keyexpantion/SB0/n3068 ), .C(\U1/keyexpantion/SB0/n3067 ), .D(
        \U1/keyexpantion/SB0/n3066 ), .E(\U1/keyexpantion/SB0/n3065 ), .F(
        \U1/keyexpantion/SB0/n3064 ), .Y(\U1/keyexpantion/SB0/n3149 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U114  ( .A0(
        \U1/keyexpantion/SB0/n3240 ), .A1(\U1/keyexpantion/SB0/n3070 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .B1(\U1/keyexpantion/SB0/n3196 ), .Y(
        \U1/keyexpantion/SB0/n3071 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U113  ( .A0(
        \U1/keyexpantion/SB0/n3122 ), .A1(\U1/keyexpantion/SB0/n3267 ), .B0(
        \U1/keyexpantion/SB0/n3072 ), .B1(\U1/keyexpantion/SB0/n3257 ), .C0(
        \U1/keyexpantion/SB0/n3071 ), .Y(\U1/keyexpantion/SB0/n3084 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U112  ( .AN(
        \U1/keyexpantion/SB0/n3076 ), .B(\U1/keyexpantion/SB0/n3075 ), .C(
        \U1/keyexpantion/SB0/n3074 ), .D(\U1/keyexpantion/SB0/n3073 ), .Y(
        \U1/keyexpantion/SB0/n3083 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U111  ( .A0(
        \U1/keyexpantion/SB0/n3260 ), .A1(\U1/keyexpantion/SB0/n3077 ), .B0(
        \U1/keyexpantion/SB0/n3251 ), .Y(\U1/keyexpantion/SB0/n3081 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U110  ( .A(
        \U1/keyexpantion/SB0/n3227 ), .B(\U1/keyexpantion/SB0/n3232 ), .Y(
        \U1/keyexpantion/SB0/n3078 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U109  ( .A0(
        \U1/keyexpantion/SB0/n3203 ), .A1(\U1/keyexpantion/SB0/n3078 ), .B0(
        \U1/keyexpantion/SB0/n3204 ), .B1(\U1/keyexpantion/SB0/n3150 ), .Y(
        \U1/keyexpantion/SB0/n3079 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U108  ( .A(
        \U1/keyexpantion/SB0/n3081 ), .B(\U1/keyexpantion/SB0/n3080 ), .C(
        \U1/keyexpantion/SB0/n3079 ), .Y(\U1/keyexpantion/SB0/n3082 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U107  ( .A(\U1/keyexpantion/SB0/n3142 ), 
        .B(\U1/keyexpantion/SB0/n3190 ), .C(\U1/keyexpantion/SB0/n3149 ), .D(
        \U1/keyexpantion/SB0/n3084 ), .E(\U1/keyexpantion/SB0/n3083 ), .F(
        \U1/keyexpantion/SB0/n3082 ), .Y(\U1/keyexpantion/SB0/n3236 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U106  ( .A(\U1/keyexpantion/SB0/n3169 ), 
        .B(\U1/keyexpantion/SB0/n3214 ), .C(\U1/keyexpantion/SB0/n3118 ), .D(
        \U1/keyexpantion/SB0/n3236 ), .Y(\U1/keyexpantion/SB0/n3098 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U105  ( .A0(
        \U1/keyexpantion/SB0/n3216 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n3085 ), .B1(\U1/keyexpantion/SB0/n3232 ), .Y(
        \U1/keyexpantion/SB0/n3086 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U104  ( .A0(
        \U1/keyexpantion/SB0/n3221 ), .A1(\U1/keyexpantion/SB0/n3239 ), .B0(
        \U1/keyexpantion/SB0/n3252 ), .B1(\U1/keyexpantion/SB0/n3260 ), .C0(
        \U1/keyexpantion/SB0/n3086 ), .Y(\U1/keyexpantion/SB0/n3097 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U103  ( .A(\U1/keyexpantion/SB0/n3087 ), 
        .Y(\U1/keyexpantion/SB0/n3090 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U102  ( .A0(
        \U1/keyexpantion/SB0/n3088 ), .A1(\U1/keyexpantion/SB0/n3193 ), .B0(
        \U1/keyexpantion/SB0/n3121 ), .B1(\U1/keyexpantion/SB0/n3173 ), .Y(
        \U1/keyexpantion/SB0/n3089 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U101  ( .A0(
        \U1/keyexpantion/SB0/n3240 ), .A1(\U1/keyexpantion/SB0/n3090 ), .B0(
        \U1/keyexpantion/SB0/n3222 ), .B1(\U1/keyexpantion/SB0/n3171 ), .C0(
        \U1/keyexpantion/SB0/n3089 ), .Y(\U1/keyexpantion/SB0/n3096 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U100  ( .A0(
        \U1/keyexpantion/SB0/n3262 ), .A1(\U1/keyexpantion/SB0/n3139 ), .B0(
        \U1/keyexpantion/SB0/n3242 ), .Y(\U1/keyexpantion/SB0/n3094 ) );
  AND4_X0P5M_A12TL \U1/keyexpantion/SB0/U99  ( .A(\U1/keyexpantion/SB0/n3094 ), 
        .B(\U1/keyexpantion/SB0/n3093 ), .C(\U1/keyexpantion/SB0/n3092 ), .D(
        \U1/keyexpantion/SB0/n3091 ), .Y(\U1/keyexpantion/SB0/n3095 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U98  ( .AN(
        \U1/keyexpantion/SB0/n3098 ), .B(\U1/keyexpantion/SB0/n3097 ), .C(
        \U1/keyexpantion/SB0/n3096 ), .D(\U1/keyexpantion/SB0/n3095 ), .Y(
        \U1/keyexpantion/ws [3]) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U97  ( .A0(
        \U1/keyexpantion/SB0/n3113 ), .A1(\U1/keyexpantion/SB0/n3228 ), .B0(
        \U1/keyexpantion/SB0/n3172 ), .Y(\U1/keyexpantion/SB0/n3110 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U96  ( .A(\U1/keyexpantion/SB0/n3101 ), .B(\U1/keyexpantion/SB0/n3100 ), .C(\U1/keyexpantion/SB0/n3099 ), .Y(
        \U1/keyexpantion/SB0/n3109 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U95  ( .A(\U1/keyexpantion/SB0/n3240 ), 
        .B(\U1/keyexpantion/SB0/n3251 ), .Y(\U1/keyexpantion/SB0/n3104 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U94  ( .A(\U1/keyexpantion/SB0/n3222 ), 
        .B(\U1/keyexpantion/SB0/n3156 ), .Y(\U1/keyexpantion/SB0/n3102 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U93  ( .A0(
        \U1/keyexpantion/SB0/n3104 ), .A1(\U1/keyexpantion/SB0/n3103 ), .B0(
        \U1/keyexpantion/SB0/n3102 ), .B1(\U1/keyexpantion/SB0/n3245 ), .C0(
        \U1/keyexpantion/SB0/n3228 ), .C1(\U1/keyexpantion/SB0/n3154 ), .Y(
        \U1/keyexpantion/SB0/n3108 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U92  ( .A0(
        \U1/keyexpantion/SB0/n3205 ), .A1(\U1/keyexpantion/SB0/n3106 ), .B0(
        \U1/keyexpantion/SB0/n3267 ), .B1(\U1/keyexpantion/SB0/n3257 ), .C0(
        \U1/keyexpantion/SB0/n3230 ), .C1(\U1/keyexpantion/SB0/n3105 ), .Y(
        \U1/keyexpantion/SB0/n3107 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U91  ( .A(\U1/keyexpantion/SB0/n3112 ), 
        .B(\U1/keyexpantion/SB0/n3111 ), .C(\U1/keyexpantion/SB0/n3110 ), .D(
        \U1/keyexpantion/SB0/n3109 ), .E(\U1/keyexpantion/SB0/n3108 ), .F(
        \U1/keyexpantion/SB0/n3107 ), .Y(\U1/keyexpantion/SB0/n3237 ) );
  AOI21_X0P5M_A12TL \U1/keyexpantion/SB0/U90  ( .A0(
        \U1/keyexpantion/SB0/n3113 ), .A1(\U1/keyexpantion/SB0/n3122 ), .B0(
        \U1/keyexpantion/SB0/n3193 ), .Y(\U1/keyexpantion/SB0/n3148 ) );
  AOI31_X0P5M_A12TL \U1/keyexpantion/SB0/U89  ( .A0(
        \U1/keyexpantion/SB0/n3217 ), .A1(\U1/keyexpantion/SB0/n3230 ), .A2(
        \U1/keyexpantion/SB0/n3170 ), .B0(\U1/keyexpantion/SB0/n3246 ), .Y(
        \U1/keyexpantion/SB0/n3147 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U88  ( .A(\U1/keyexpantion/SB0/n3117 ), .B(\U1/keyexpantion/SB0/n3116 ), .C(\U1/keyexpantion/SB0/n3115 ), .D(
        \U1/keyexpantion/SB0/n3114 ), .Y(\U1/keyexpantion/SB0/n3144 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U87  ( .A(\U1/keyexpantion/SB0/n3118 ), 
        .Y(\U1/keyexpantion/SB0/n3141 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U86  ( .A(\U1/keyexpantion/SB0/n3119 ), 
        .Y(\U1/keyexpantion/SB0/n3135 ) );
  OAI21B_X0P5M_A12TL \U1/keyexpantion/SB0/U85  ( .A0(
        \U1/keyexpantion/SB0/n3121 ), .A1(\U1/keyexpantion/SB0/n3258 ), .B0N(
        \U1/keyexpantion/SB0/n3120 ), .Y(\U1/keyexpantion/SB0/n3134 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U84  ( .A0(
        \U1/keyexpantion/SB0/n3265 ), .A1(\U1/keyexpantion/SB0/n3122 ), .B0(
        \U1/keyexpantion/SB0/n3172 ), .B1(\U1/keyexpantion/SB0/n3232 ), .C0(
        \U1/keyexpantion/SB0/n3246 ), .C1(\U1/keyexpantion/SB0/n3267 ), .Y(
        \U1/keyexpantion/SB0/n3133 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U83  ( .AN(
        \U1/keyexpantion/SB0/n3126 ), .B(\U1/keyexpantion/SB0/n3125 ), .C(
        \U1/keyexpantion/SB0/n3124 ), .D(\U1/keyexpantion/SB0/n3123 ), .Y(
        \U1/keyexpantion/SB0/n3132 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U82  ( .A(\U1/keyexpantion/SB0/n3130 ), .B(\U1/keyexpantion/SB0/n3129 ), .C(\U1/keyexpantion/SB0/n3128 ), .D(
        \U1/keyexpantion/SB0/n3127 ), .Y(\U1/keyexpantion/SB0/n3131 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U81  ( .A(\U1/keyexpantion/SB0/n3136 ), 
        .B(\U1/keyexpantion/SB0/n3135 ), .C(\U1/keyexpantion/SB0/n3134 ), .D(
        \U1/keyexpantion/SB0/n3133 ), .E(\U1/keyexpantion/SB0/n3132 ), .F(
        \U1/keyexpantion/SB0/n3131 ), .Y(\U1/keyexpantion/SB0/n3137 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U80  ( .A(\U1/keyexpantion/SB0/n3137 ), 
        .Y(\U1/keyexpantion/SB0/n3215 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U79  ( .A0(
        \U1/keyexpantion/SB0/n3205 ), .A1(\U1/keyexpantion/SB0/n3227 ), .B0(
        \U1/keyexpantion/SB0/n3267 ), .B1(\U1/keyexpantion/SB0/n3266 ), .Y(
        \U1/keyexpantion/SB0/n3138 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U78  ( .A0(
        \U1/keyexpantion/SB0/n3195 ), .A1(\U1/keyexpantion/SB0/n3139 ), .B0(
        \U1/keyexpantion/SB0/n3219 ), .B1(\U1/keyexpantion/SB0/n3241 ), .C0(
        \U1/keyexpantion/SB0/n3138 ), .Y(\U1/keyexpantion/SB0/n3140 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U77  ( .AN(
        \U1/keyexpantion/SB0/n3142 ), .B(\U1/keyexpantion/SB0/n3141 ), .C(
        \U1/keyexpantion/SB0/n3215 ), .D(\U1/keyexpantion/SB0/n3140 ), .Y(
        \U1/keyexpantion/SB0/n3143 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U76  ( .A(\U1/keyexpantion/SB0/n3148 ), 
        .B(\U1/keyexpantion/SB0/n3147 ), .C(\U1/keyexpantion/SB0/n3146 ), .D(
        \U1/keyexpantion/SB0/n3145 ), .E(\U1/keyexpantion/SB0/n3144 ), .F(
        \U1/keyexpantion/SB0/n3143 ), .Y(\U1/keyexpantion/SB0/n3213 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U75  ( .A(\U1/keyexpantion/SB0/n3149 ), 
        .Y(\U1/keyexpantion/SB0/n3153 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U74  ( .A0(
        \U1/keyexpantion/SB0/n3151 ), .A1(\U1/keyexpantion/SB0/n3150 ), .B0(
        \U1/keyexpantion/SB0/n3197 ), .B1(\U1/keyexpantion/SB0/n3156 ), .Y(
        \U1/keyexpantion/SB0/n3152 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U73  ( .A0(
        \U1/keyexpantion/SB0/n3246 ), .A1(\U1/keyexpantion/SB0/n3154 ), .B0(
        \U1/keyexpantion/SB0/n3153 ), .C0(\U1/keyexpantion/SB0/n3152 ), .Y(
        \U1/keyexpantion/SB0/n3168 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U72  ( .A0(
        \U1/keyexpantion/SB0/n3155 ), .A1(\U1/keyexpantion/SB0/n3218 ), .B0(
        \U1/keyexpantion/SB0/n3247 ), .Y(\U1/keyexpantion/SB0/n3160 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U71  ( .A0(
        \U1/keyexpantion/SB0/n3156 ), .A1(\U1/keyexpantion/SB0/n3221 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n3159 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U70  ( .A(\U1/keyexpantion/SB0/n3160 ), .B(\U1/keyexpantion/SB0/n3159 ), .C(\U1/keyexpantion/SB0/n3158 ), .D(
        \U1/keyexpantion/SB0/n3157 ), .Y(\U1/keyexpantion/SB0/n3167 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U69  ( .A(\U1/keyexpantion/SB0/n3198 ), 
        .B(\U1/keyexpantion/SB0/n3161 ), .Y(\U1/keyexpantion/SB0/n3165 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U68  ( .A(\U1/keyexpantion/SB0/n3162 ), 
        .B(\U1/keyexpantion/SB0/n3203 ), .Y(\U1/keyexpantion/SB0/n3164 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U67  ( .A0(
        \U1/keyexpantion/SB0/n3165 ), .A1(\U1/keyexpantion/SB0/n3264 ), .B0(
        \U1/keyexpantion/SB0/n3164 ), .B1(\U1/keyexpantion/SB0/n3228 ), .C0(
        \U1/keyexpantion/SB0/n3163 ), .C1(\U1/keyexpantion/SB0/n3229 ), .Y(
        \U1/keyexpantion/SB0/n3166 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U66  ( .A(\U1/keyexpantion/SB0/n3237 ), 
        .B(\U1/keyexpantion/SB0/n3213 ), .C(\U1/keyexpantion/SB0/n3169 ), .D(
        \U1/keyexpantion/SB0/n3168 ), .E(\U1/keyexpantion/SB0/n3167 ), .F(
        \U1/keyexpantion/SB0/n3166 ), .Y(\U1/keyexpantion/ws [4]) );
  AOI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U65  ( .A1N(
        \U1/keyexpantion/SB0/n3171 ), .A0(\U1/keyexpantion/SB0/n3170 ), .B0(
        \U1/keyexpantion/SB0/n3227 ), .Y(\U1/keyexpantion/SB0/n3187 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U64  ( .A(\U1/keyexpantion/SB0/n3240 ), 
        .B(\U1/keyexpantion/SB0/n3221 ), .Y(\U1/keyexpantion/SB0/n3174 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U63  ( .A0(
        \U1/keyexpantion/SB0/n3264 ), .A1(\U1/keyexpantion/SB0/n3175 ), .B0(
        \U1/keyexpantion/SB0/n3174 ), .B1(\U1/keyexpantion/SB0/n3267 ), .C0(
        \U1/keyexpantion/SB0/n3173 ), .C1(\U1/keyexpantion/SB0/n3172 ), .Y(
        \U1/keyexpantion/SB0/n3186 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U62  ( .A(\U1/keyexpantion/SB0/n3176 ), 
        .Y(\U1/keyexpantion/SB0/n3179 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U61  ( .AN(
        \U1/keyexpantion/SB0/n3180 ), .B(\U1/keyexpantion/SB0/n3179 ), .C(
        \U1/keyexpantion/SB0/n3178 ), .D(\U1/keyexpantion/SB0/n3177 ), .Y(
        \U1/keyexpantion/SB0/n3185 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U60  ( .A(\U1/keyexpantion/SB0/n3183 ), .B(\U1/keyexpantion/SB0/n3182 ), .C(\U1/keyexpantion/SB0/n3181 ), .Y(
        \U1/keyexpantion/SB0/n3184 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U59  ( .A(\U1/keyexpantion/SB0/n3189 ), 
        .B(\U1/keyexpantion/SB0/n3188 ), .C(\U1/keyexpantion/SB0/n3187 ), .D(
        \U1/keyexpantion/SB0/n3186 ), .E(\U1/keyexpantion/SB0/n3185 ), .F(
        \U1/keyexpantion/SB0/n3184 ), .Y(\U1/keyexpantion/SB0/n3238 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U58  ( .A(\U1/keyexpantion/SB0/n3190 ), 
        .Y(\U1/keyexpantion/SB0/n3192 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U57  ( .A0(
        \U1/keyexpantion/SB0/n3251 ), .A1(\U1/keyexpantion/SB0/n3248 ), .B0(
        \U1/keyexpantion/SB0/n3252 ), .B1(\U1/keyexpantion/SB0/n3250 ), .Y(
        \U1/keyexpantion/SB0/n3191 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U56  ( .A0(
        \U1/keyexpantion/SB0/n3227 ), .A1(\U1/keyexpantion/SB0/n3193 ), .B0(
        \U1/keyexpantion/SB0/n3192 ), .C0(\U1/keyexpantion/SB0/n3191 ), .Y(
        \U1/keyexpantion/SB0/n3212 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U55  ( .A0(
        \U1/keyexpantion/SB0/n3195 ), .A1(\U1/keyexpantion/SB0/n3251 ), .B0(
        \U1/keyexpantion/SB0/n3194 ), .Y(\U1/keyexpantion/SB0/n3201 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U54  ( .A0(
        \U1/keyexpantion/SB0/n3198 ), .A1(\U1/keyexpantion/SB0/n3197 ), .B0(
        \U1/keyexpantion/SB0/n3196 ), .Y(\U1/keyexpantion/SB0/n3200 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U53  ( .AN(
        \U1/keyexpantion/SB0/n3202 ), .B(\U1/keyexpantion/SB0/n3201 ), .C(
        \U1/keyexpantion/SB0/n3200 ), .D(\U1/keyexpantion/SB0/n3199 ), .Y(
        \U1/keyexpantion/SB0/n3211 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U52  ( .A0(
        \U1/keyexpantion/SB0/n3247 ), .A1(\U1/keyexpantion/SB0/n3204 ), .B0(
        \U1/keyexpantion/SB0/n3203 ), .Y(\U1/keyexpantion/SB0/n3208 ) );
  OA22_X0P5M_A12TL \U1/keyexpantion/SB0/U51  ( .A0(\U1/keyexpantion/SB0/n3229 ), .A1(\U1/keyexpantion/SB0/n3206 ), .B0(\U1/keyexpantion/SB0/n3266 ), .B1(
        \U1/keyexpantion/SB0/n3205 ), .Y(\U1/keyexpantion/SB0/n3207 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U50  ( .A0(
        \U1/keyexpantion/SB0/n3209 ), .A1(\U1/keyexpantion/SB0/n3228 ), .B0(
        \U1/keyexpantion/SB0/n3208 ), .C0(\U1/keyexpantion/SB0/n3207 ), .Y(
        \U1/keyexpantion/SB0/n3210 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U49  ( .A(\U1/keyexpantion/SB0/n3238 ), 
        .B(\U1/keyexpantion/SB0/n3214 ), .C(\U1/keyexpantion/SB0/n3213 ), .D(
        \U1/keyexpantion/SB0/n3212 ), .E(\U1/keyexpantion/SB0/n3211 ), .F(
        \U1/keyexpantion/SB0/n3210 ), .Y(\U1/keyexpantion/ws [5]) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U48  ( .A0(
        \U1/keyexpantion/SB0/n3217 ), .A1(\U1/keyexpantion/SB0/n3257 ), .B0(
        \U1/keyexpantion/SB0/n3216 ), .B1(\U1/keyexpantion/SB0/n3264 ), .C0(
        \U1/keyexpantion/SB0/n3215 ), .Y(\U1/keyexpantion/SB0/n3235 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U47  ( .A0(
        \U1/keyexpantion/SB0/n3218 ), .A1(\U1/keyexpantion/SB0/n3262 ), .B0(
        \U1/keyexpantion/SB0/n3251 ), .Y(\U1/keyexpantion/SB0/n3226 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U46  ( .A0(
        \U1/keyexpantion/SB0/n3242 ), .A1(\U1/keyexpantion/SB0/n3219 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n3225 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U45  ( .A0(
        \U1/keyexpantion/SB0/n3222 ), .A1(\U1/keyexpantion/SB0/n3221 ), .B0(
        \U1/keyexpantion/SB0/n3220 ), .Y(\U1/keyexpantion/SB0/n3224 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U44  ( .A(\U1/keyexpantion/SB0/n3226 ), .B(\U1/keyexpantion/SB0/n3225 ), .C(\U1/keyexpantion/SB0/n3224 ), .D(
        \U1/keyexpantion/SB0/n3223 ), .Y(\U1/keyexpantion/SB0/n3234 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U43  ( .A(\U1/keyexpantion/SB0/n3257 ), .B(\U1/keyexpantion/SB0/n3227 ), .Y(\U1/keyexpantion/SB0/n3259 ) );
  NOR2_X0P5A_A12TL \U1/keyexpantion/SB0/U42  ( .A(\U1/keyexpantion/SB0/n3247 ), 
        .B(\U1/keyexpantion/SB0/n3259 ), .Y(\U1/keyexpantion/SB0/n3231 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U41  ( .A0(
        \U1/keyexpantion/SB0/n3245 ), .A1(\U1/keyexpantion/SB0/n3232 ), .B0(
        \U1/keyexpantion/SB0/n3231 ), .B1(\U1/keyexpantion/SB0/n3230 ), .C0(
        \U1/keyexpantion/SB0/n3229 ), .C1(\U1/keyexpantion/SB0/n3228 ), .Y(
        \U1/keyexpantion/SB0/n3233 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U40  ( .A(\U1/keyexpantion/SB0/n3238 ), 
        .B(\U1/keyexpantion/SB0/n3237 ), .C(\U1/keyexpantion/SB0/n3236 ), .D(
        \U1/keyexpantion/SB0/n3235 ), .E(\U1/keyexpantion/SB0/n3234 ), .F(
        \U1/keyexpantion/SB0/n3233 ), .Y(\U1/keyexpantion/ws [6]) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U39  ( .A0(
        \U1/keyexpantion/SB0/n3242 ), .A1(\U1/keyexpantion/SB0/n3241 ), .B0(
        \U1/keyexpantion/SB0/n3240 ), .B1(\U1/keyexpantion/SB0/n3239 ), .Y(
        \U1/keyexpantion/SB0/n3243 ) );
  OAI211_X0P5M_A12TL \U1/keyexpantion/SB0/U38  ( .A0(
        \U1/keyexpantion/SB0/n3246 ), .A1(\U1/keyexpantion/SB0/n3245 ), .B0(
        \U1/keyexpantion/SB0/n3244 ), .C0(\U1/keyexpantion/SB0/n3243 ), .Y(
        \U1/keyexpantion/SB0/n3270 ) );
  OAI2XB1_X0P5M_A12TL \U1/keyexpantion/SB0/U37  ( .A1N(
        \U1/keyexpantion/SB0/n3249 ), .A0(\U1/keyexpantion/SB0/n3248 ), .B0(
        \U1/keyexpantion/SB0/n3247 ), .Y(\U1/keyexpantion/SB0/n3256 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U36  ( .A0(
        \U1/keyexpantion/SB0/n3252 ), .A1(\U1/keyexpantion/SB0/n3251 ), .B0(
        \U1/keyexpantion/SB0/n3250 ), .Y(\U1/keyexpantion/SB0/n3255 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U35  ( .A(\U1/keyexpantion/SB0/n3256 ), .B(\U1/keyexpantion/SB0/n3255 ), .C(\U1/keyexpantion/SB0/n3254 ), .D(
        \U1/keyexpantion/SB0/n3253 ), .Y(\U1/keyexpantion/SB0/n3269 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U34  ( .A(\U1/keyexpantion/SB0/n3258 ), .B(\U1/keyexpantion/SB0/n3257 ), .Y(\U1/keyexpantion/SB0/n3261 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U33  ( .A0(
        \U1/keyexpantion/SB0/n3262 ), .A1(\U1/keyexpantion/SB0/n3261 ), .B0(
        \U1/keyexpantion/SB0/n3260 ), .B1(\U1/keyexpantion/SB0/n3259 ), .Y(
        \U1/keyexpantion/SB0/n3263 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U32  ( .A0(
        \U1/keyexpantion/SB0/n3267 ), .A1(\U1/keyexpantion/SB0/n3266 ), .B0(
        \U1/keyexpantion/SB0/n3265 ), .B1(\U1/keyexpantion/SB0/n3264 ), .C0(
        \U1/keyexpantion/SB0/n3263 ), .Y(\U1/keyexpantion/SB0/n3268 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U31  ( .A(\U1/keyexpantion/SB0/n3273 ), 
        .B(\U1/keyexpantion/SB0/n3272 ), .C(\U1/keyexpantion/SB0/n3271 ), .D(
        \U1/keyexpantion/SB0/n3270 ), .E(\U1/keyexpantion/SB0/n3269 ), .F(
        \U1/keyexpantion/SB0/n3268 ), .Y(\U1/keyexpantion/ws [7]) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U30  ( .A(\U1/keyexpantion/SB0/n3276 ), .B(\U1/keyexpantion/SB0/n3275 ), .C(\U1/keyexpantion/SB0/n3274 ), .Y(
        \U1/keyexpantion/SB0/n3299 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U29  ( .A0(
        \U1/keyexpantion/SB0/n3277 ), .A1(\U1/keyexpantion/SB0/n3333 ), .B0(
        \U1/keyexpantion/SB0/n3349 ), .Y(\U1/keyexpantion/SB0/n3282 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U28  ( .A0(
        \U1/keyexpantion/SB0/n3342 ), .A1(\U1/keyexpantion/SB0/n3279 ), .B0(
        \U1/keyexpantion/SB0/n3278 ), .B1(\U1/keyexpantion/SB0/n3343 ), .Y(
        \U1/keyexpantion/SB0/n3280 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U27  ( .A(\U1/keyexpantion/SB0/n3282 ), .B(\U1/keyexpantion/SB0/n3281 ), .C(\U1/keyexpantion/SB0/n3280 ), .Y(
        \U1/keyexpantion/SB0/n3298 ) );
  AOI22_X0P5M_A12TL \U1/keyexpantion/SB0/U26  ( .A0(
        \U1/keyexpantion/SB0/n3285 ), .A1(\U1/keyexpantion/SB0/n3308 ), .B0(
        \U1/keyexpantion/SB0/n3284 ), .B1(\U1/keyexpantion/SB0/n3283 ), .Y(
        \U1/keyexpantion/SB0/n3286 ) );
  OAI221_X0P5M_A12TL \U1/keyexpantion/SB0/U25  ( .A0(
        \U1/keyexpantion/SB0/n3290 ), .A1(\U1/keyexpantion/SB0/n3289 ), .B0(
        \U1/keyexpantion/SB0/n3288 ), .B1(\U1/keyexpantion/SB0/n3287 ), .C0(
        \U1/keyexpantion/SB0/n3286 ), .Y(\U1/keyexpantion/SB0/n3297 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U24  ( .A(\U1/keyexpantion/SB0/n3338 ), .B(\U1/keyexpantion/SB0/n3291 ), .Y(\U1/keyexpantion/SB0/n3292 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U23  ( .AN(
        \U1/keyexpantion/SB0/n3295 ), .B(\U1/keyexpantion/SB0/n3294 ), .C(
        \U1/keyexpantion/SB0/n3293 ), .D(\U1/keyexpantion/SB0/n3292 ), .Y(
        \U1/keyexpantion/SB0/n3296 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U22  ( .A(\U1/keyexpantion/SB0/n3301 ), 
        .B(\U1/keyexpantion/SB0/n3300 ), .C(\U1/keyexpantion/SB0/n3299 ), .D(
        \U1/keyexpantion/SB0/n3298 ), .E(\U1/keyexpantion/SB0/n3297 ), .F(
        \U1/keyexpantion/SB0/n3296 ), .Y(\U1/keyexpantion/SB0/n3360 ) );
  OR4_X0P5M_A12TL \U1/keyexpantion/SB0/U21  ( .A(\U1/keyexpantion/SB0/n3304 ), 
        .B(\U1/keyexpantion/SB0/n3303 ), .C(\U1/keyexpantion/SB0/n3302 ), .D(
        \U1/keyexpantion/SB0/n3360 ), .Y(\U1/keyexpantion/SB0/n3329 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U20  ( .A0(
        \U1/keyexpantion/SB0/n3306 ), .A1(\U1/keyexpantion/SB0/n3317 ), .B0(
        \U1/keyexpantion/SB0/n3353 ), .B1(\U1/keyexpantion/SB0/n3305 ), .Y(
        \U1/keyexpantion/SB0/n3307 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U19  ( .A0(
        \U1/keyexpantion/SB0/n3331 ), .A1(\U1/keyexpantion/SB0/n3343 ), .B0(
        \U1/keyexpantion/SB0/n3334 ), .B1(\U1/keyexpantion/SB0/n3308 ), .C0(
        \U1/keyexpantion/SB0/n3307 ), .Y(\U1/keyexpantion/SB0/n3328 ) );
  OAI22_X0P5M_A12TL \U1/keyexpantion/SB0/U18  ( .A0(
        \U1/keyexpantion/SB0/n3312 ), .A1(\U1/keyexpantion/SB0/n3311 ), .B0(
        \U1/keyexpantion/SB0/n3310 ), .B1(\U1/keyexpantion/SB0/n3309 ), .Y(
        \U1/keyexpantion/SB0/n3313 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U17  ( .A0(
        \U1/keyexpantion/SB0/n3316 ), .A1(\U1/keyexpantion/SB0/n3315 ), .B0(
        \U1/keyexpantion/SB0/n3314 ), .B1(\U1/keyexpantion/SB0/n3339 ), .C0(
        \U1/keyexpantion/SB0/n3313 ), .Y(\U1/keyexpantion/SB0/n3327 ) );
  NAND2_X0P5A_A12TL \U1/keyexpantion/SB0/U16  ( .A(\U1/keyexpantion/SB0/n3318 ), .B(\U1/keyexpantion/SB0/n3317 ), .Y(\U1/keyexpantion/SB0/n3325 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U15  ( .A(\U1/keyexpantion/SB0/n3319 ), 
        .Y(\U1/keyexpantion/SB0/n3324 ) );
  NAND3_X0P5A_A12TL \U1/keyexpantion/SB0/U14  ( .A(\U1/keyexpantion/SB0/n3322 ), .B(\U1/keyexpantion/SB0/n3321 ), .C(\U1/keyexpantion/SB0/n3320 ), .Y(
        \U1/keyexpantion/SB0/n3323 ) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U13  ( .A0(
        \U1/keyexpantion/SB0/n3340 ), .A1(\U1/keyexpantion/SB0/n3325 ), .B0(
        \U1/keyexpantion/SB0/n3332 ), .B1(\U1/keyexpantion/SB0/n3324 ), .C0(
        \U1/keyexpantion/SB0/n3323 ), .Y(\U1/keyexpantion/SB0/n3326 ) );
  NAND4B_X0P5M_A12TL \U1/keyexpantion/SB0/U12  ( .AN(
        \U1/keyexpantion/SB0/n3329 ), .B(\U1/keyexpantion/SB0/n3328 ), .C(
        \U1/keyexpantion/SB0/n3327 ), .D(\U1/keyexpantion/SB0/n3326 ), .Y(
        \U1/keyexpantion/ws [8]) );
  AOI221_X0P5M_A12TL \U1/keyexpantion/SB0/U11  ( .A0(
        \U1/keyexpantion/SB0/n3334 ), .A1(\U1/keyexpantion/SB0/n3333 ), .B0(
        \U1/keyexpantion/SB0/n3332 ), .B1(\U1/keyexpantion/SB0/n3331 ), .C0(
        \U1/keyexpantion/SB0/n3330 ), .Y(\U1/keyexpantion/SB0/n3335 ) );
  INV_X0P5B_A12TL \U1/keyexpantion/SB0/U10  ( .A(\U1/keyexpantion/SB0/n3335 ), 
        .Y(\U1/keyexpantion/SB0/n3359 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U9  ( .A0(\U1/keyexpantion/SB0/n3348 ), .A1(\U1/keyexpantion/SB0/n3337 ), .B0(\U1/keyexpantion/SB0/n3336 ), .Y(
        \U1/keyexpantion/SB0/n3347 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U8  ( .A0(\U1/keyexpantion/SB0/n3340 ), .A1(\U1/keyexpantion/SB0/n3339 ), .B0(\U1/keyexpantion/SB0/n3338 ), .Y(
        \U1/keyexpantion/SB0/n3346 ) );
  OAI21_X0P5M_A12TL \U1/keyexpantion/SB0/U7  ( .A0(\U1/keyexpantion/SB0/n3343 ), .A1(\U1/keyexpantion/SB0/n3342 ), .B0(\U1/keyexpantion/SB0/n3341 ), .Y(
        \U1/keyexpantion/SB0/n3345 ) );
  NAND4_X0P5A_A12TL \U1/keyexpantion/SB0/U6  ( .A(\U1/keyexpantion/SB0/n3347 ), 
        .B(\U1/keyexpantion/SB0/n3346 ), .C(\U1/keyexpantion/SB0/n3345 ), .D(
        \U1/keyexpantion/SB0/n3344 ), .Y(\U1/keyexpantion/SB0/n3358 ) );
  NOR3_X0P5A_A12TL \U1/keyexpantion/SB0/U5  ( .A(\U1/keyexpantion/SB0/n3350 ), 
        .B(\U1/keyexpantion/SB0/n3349 ), .C(\U1/keyexpantion/SB0/n3348 ), .Y(
        \U1/keyexpantion/SB0/n3354 ) );
  OAI222_X0P5M_A12TL \U1/keyexpantion/SB0/U4  ( .A0(
        \U1/keyexpantion/SB0/n3356 ), .A1(\U1/keyexpantion/SB0/n3355 ), .B0(
        \U1/keyexpantion/SB0/n3354 ), .B1(\U1/keyexpantion/SB0/n3353 ), .C0(
        \U1/keyexpantion/SB0/n3352 ), .C1(\U1/keyexpantion/SB0/n3351 ), .Y(
        \U1/keyexpantion/SB0/n3357 ) );
  OR6_X0P5M_A12TL \U1/keyexpantion/SB0/U3  ( .A(\U1/keyexpantion/SB0/n3362 ), 
        .B(\U1/keyexpantion/SB0/n3361 ), .C(\U1/keyexpantion/SB0/n3360 ), .D(
        \U1/keyexpantion/SB0/n3359 ), .E(\U1/keyexpantion/SB0/n3358 ), .F(
        \U1/keyexpantion/SB0/n3357 ), .Y(\U1/keyexpantion/ws [9]) );
endmodule

